magic
tech sky130A
magscale 1 2
timestamp 1644999282
<< obsli1 >>
rect 1104 2159 197311 198033
<< obsm1 >>
rect 1104 620 197786 198348
<< metal2 >>
rect 570 199504 626 200304
rect 1766 199504 1822 200304
rect 2962 199504 3018 200304
rect 4158 199504 4214 200304
rect 5354 199504 5410 200304
rect 6550 199504 6606 200304
rect 7746 199504 7802 200304
rect 8942 199504 8998 200304
rect 10230 199504 10286 200304
rect 11426 199504 11482 200304
rect 12622 199504 12678 200304
rect 13818 199504 13874 200304
rect 15014 199504 15070 200304
rect 16210 199504 16266 200304
rect 17406 199504 17462 200304
rect 18694 199504 18750 200304
rect 19890 199504 19946 200304
rect 21086 199504 21142 200304
rect 22282 199504 22338 200304
rect 23478 199504 23534 200304
rect 24674 199504 24730 200304
rect 25870 199504 25926 200304
rect 27066 199504 27122 200304
rect 28354 199504 28410 200304
rect 29550 199504 29606 200304
rect 30746 199504 30802 200304
rect 31942 199504 31998 200304
rect 33138 199504 33194 200304
rect 34334 199504 34390 200304
rect 35530 199504 35586 200304
rect 36818 199504 36874 200304
rect 38014 199504 38070 200304
rect 39210 199504 39266 200304
rect 40406 199504 40462 200304
rect 41602 199504 41658 200304
rect 42798 199504 42854 200304
rect 43994 199504 44050 200304
rect 45190 199504 45246 200304
rect 46478 199504 46534 200304
rect 47674 199504 47730 200304
rect 48870 199504 48926 200304
rect 50066 199504 50122 200304
rect 51262 199504 51318 200304
rect 52458 199504 52514 200304
rect 53654 199504 53710 200304
rect 54942 199504 54998 200304
rect 56138 199504 56194 200304
rect 57334 199504 57390 200304
rect 58530 199504 58586 200304
rect 59726 199504 59782 200304
rect 60922 199504 60978 200304
rect 62118 199504 62174 200304
rect 63314 199504 63370 200304
rect 64602 199504 64658 200304
rect 65798 199504 65854 200304
rect 66994 199504 67050 200304
rect 68190 199504 68246 200304
rect 69386 199504 69442 200304
rect 70582 199504 70638 200304
rect 71778 199504 71834 200304
rect 73066 199504 73122 200304
rect 74262 199504 74318 200304
rect 75458 199504 75514 200304
rect 76654 199504 76710 200304
rect 77850 199504 77906 200304
rect 79046 199504 79102 200304
rect 80242 199504 80298 200304
rect 81438 199504 81494 200304
rect 82726 199504 82782 200304
rect 83922 199504 83978 200304
rect 85118 199504 85174 200304
rect 86314 199504 86370 200304
rect 87510 199504 87566 200304
rect 88706 199504 88762 200304
rect 89902 199504 89958 200304
rect 91190 199504 91246 200304
rect 92386 199504 92442 200304
rect 93582 199504 93638 200304
rect 94778 199504 94834 200304
rect 95974 199504 96030 200304
rect 97170 199504 97226 200304
rect 98366 199504 98422 200304
rect 99654 199504 99710 200304
rect 100850 199504 100906 200304
rect 102046 199504 102102 200304
rect 103242 199504 103298 200304
rect 104438 199504 104494 200304
rect 105634 199504 105690 200304
rect 106830 199504 106886 200304
rect 108026 199504 108082 200304
rect 109314 199504 109370 200304
rect 110510 199504 110566 200304
rect 111706 199504 111762 200304
rect 112902 199504 112958 200304
rect 114098 199504 114154 200304
rect 115294 199504 115350 200304
rect 116490 199504 116546 200304
rect 117778 199504 117834 200304
rect 118974 199504 119030 200304
rect 120170 199504 120226 200304
rect 121366 199504 121422 200304
rect 122562 199504 122618 200304
rect 123758 199504 123814 200304
rect 124954 199504 125010 200304
rect 126150 199504 126206 200304
rect 127438 199504 127494 200304
rect 128634 199504 128690 200304
rect 129830 199504 129886 200304
rect 131026 199504 131082 200304
rect 132222 199504 132278 200304
rect 133418 199504 133474 200304
rect 134614 199504 134670 200304
rect 135902 199504 135958 200304
rect 137098 199504 137154 200304
rect 138294 199504 138350 200304
rect 139490 199504 139546 200304
rect 140686 199504 140742 200304
rect 141882 199504 141938 200304
rect 143078 199504 143134 200304
rect 144274 199504 144330 200304
rect 145562 199504 145618 200304
rect 146758 199504 146814 200304
rect 147954 199504 148010 200304
rect 149150 199504 149206 200304
rect 150346 199504 150402 200304
rect 151542 199504 151598 200304
rect 152738 199504 152794 200304
rect 154026 199504 154082 200304
rect 155222 199504 155278 200304
rect 156418 199504 156474 200304
rect 157614 199504 157670 200304
rect 158810 199504 158866 200304
rect 160006 199504 160062 200304
rect 161202 199504 161258 200304
rect 162398 199504 162454 200304
rect 163686 199504 163742 200304
rect 164882 199504 164938 200304
rect 166078 199504 166134 200304
rect 167274 199504 167330 200304
rect 168470 199504 168526 200304
rect 169666 199504 169722 200304
rect 170862 199504 170918 200304
rect 172150 199504 172206 200304
rect 173346 199504 173402 200304
rect 174542 199504 174598 200304
rect 175738 199504 175794 200304
rect 176934 199504 176990 200304
rect 178130 199504 178186 200304
rect 179326 199504 179382 200304
rect 180522 199504 180578 200304
rect 181810 199504 181866 200304
rect 183006 199504 183062 200304
rect 184202 199504 184258 200304
rect 185398 199504 185454 200304
rect 186594 199504 186650 200304
rect 187790 199504 187846 200304
rect 188986 199504 189042 200304
rect 190274 199504 190330 200304
rect 191470 199504 191526 200304
rect 192666 199504 192722 200304
rect 193862 199504 193918 200304
rect 195058 199504 195114 200304
rect 196254 199504 196310 200304
rect 197450 199504 197506 200304
rect 662 0 718 800
rect 2042 0 2098 800
rect 3422 0 3478 800
rect 4802 0 4858 800
rect 6182 0 6238 800
rect 7562 0 7618 800
rect 8942 0 8998 800
rect 10322 0 10378 800
rect 11702 0 11758 800
rect 13082 0 13138 800
rect 14462 0 14518 800
rect 15842 0 15898 800
rect 17222 0 17278 800
rect 18602 0 18658 800
rect 19982 0 20038 800
rect 21362 0 21418 800
rect 22834 0 22890 800
rect 24214 0 24270 800
rect 25594 0 25650 800
rect 26974 0 27030 800
rect 28354 0 28410 800
rect 29734 0 29790 800
rect 31114 0 31170 800
rect 32494 0 32550 800
rect 33874 0 33930 800
rect 35254 0 35310 800
rect 36634 0 36690 800
rect 38014 0 38070 800
rect 39394 0 39450 800
rect 40774 0 40830 800
rect 42154 0 42210 800
rect 43534 0 43590 800
rect 45006 0 45062 800
rect 46386 0 46442 800
rect 47766 0 47822 800
rect 49146 0 49202 800
rect 50526 0 50582 800
rect 51906 0 51962 800
rect 53286 0 53342 800
rect 54666 0 54722 800
rect 56046 0 56102 800
rect 57426 0 57482 800
rect 58806 0 58862 800
rect 60186 0 60242 800
rect 61566 0 61622 800
rect 62946 0 63002 800
rect 64326 0 64382 800
rect 65706 0 65762 800
rect 67178 0 67234 800
rect 68558 0 68614 800
rect 69938 0 69994 800
rect 71318 0 71374 800
rect 72698 0 72754 800
rect 74078 0 74134 800
rect 75458 0 75514 800
rect 76838 0 76894 800
rect 78218 0 78274 800
rect 79598 0 79654 800
rect 80978 0 81034 800
rect 82358 0 82414 800
rect 83738 0 83794 800
rect 85118 0 85174 800
rect 86498 0 86554 800
rect 87878 0 87934 800
rect 89350 0 89406 800
rect 90730 0 90786 800
rect 92110 0 92166 800
rect 93490 0 93546 800
rect 94870 0 94926 800
rect 96250 0 96306 800
rect 97630 0 97686 800
rect 99010 0 99066 800
rect 100390 0 100446 800
rect 101770 0 101826 800
rect 103150 0 103206 800
rect 104530 0 104586 800
rect 105910 0 105966 800
rect 107290 0 107346 800
rect 108670 0 108726 800
rect 110050 0 110106 800
rect 111522 0 111578 800
rect 112902 0 112958 800
rect 114282 0 114338 800
rect 115662 0 115718 800
rect 117042 0 117098 800
rect 118422 0 118478 800
rect 119802 0 119858 800
rect 121182 0 121238 800
rect 122562 0 122618 800
rect 123942 0 123998 800
rect 125322 0 125378 800
rect 126702 0 126758 800
rect 128082 0 128138 800
rect 129462 0 129518 800
rect 130842 0 130898 800
rect 132222 0 132278 800
rect 133694 0 133750 800
rect 135074 0 135130 800
rect 136454 0 136510 800
rect 137834 0 137890 800
rect 139214 0 139270 800
rect 140594 0 140650 800
rect 141974 0 142030 800
rect 143354 0 143410 800
rect 144734 0 144790 800
rect 146114 0 146170 800
rect 147494 0 147550 800
rect 148874 0 148930 800
rect 150254 0 150310 800
rect 151634 0 151690 800
rect 153014 0 153070 800
rect 154394 0 154450 800
rect 155866 0 155922 800
rect 157246 0 157302 800
rect 158626 0 158682 800
rect 160006 0 160062 800
rect 161386 0 161442 800
rect 162766 0 162822 800
rect 164146 0 164202 800
rect 165526 0 165582 800
rect 166906 0 166962 800
rect 168286 0 168342 800
rect 169666 0 169722 800
rect 171046 0 171102 800
rect 172426 0 172482 800
rect 173806 0 173862 800
rect 175186 0 175242 800
rect 176566 0 176622 800
rect 178038 0 178094 800
rect 179418 0 179474 800
rect 180798 0 180854 800
rect 182178 0 182234 800
rect 183558 0 183614 800
rect 184938 0 184994 800
rect 186318 0 186374 800
rect 187698 0 187754 800
rect 189078 0 189134 800
rect 190458 0 190514 800
rect 191838 0 191894 800
rect 193218 0 193274 800
rect 194598 0 194654 800
rect 195978 0 196034 800
rect 197358 0 197414 800
<< obsm2 >>
rect 18 199448 514 199594
rect 682 199448 1710 199594
rect 1878 199448 2906 199594
rect 3074 199448 4102 199594
rect 4270 199448 5298 199594
rect 5466 199448 6494 199594
rect 6662 199448 7690 199594
rect 7858 199448 8886 199594
rect 9054 199448 10174 199594
rect 10342 199448 11370 199594
rect 11538 199448 12566 199594
rect 12734 199448 13762 199594
rect 13930 199448 14958 199594
rect 15126 199448 16154 199594
rect 16322 199448 17350 199594
rect 17518 199448 18638 199594
rect 18806 199448 19834 199594
rect 20002 199448 21030 199594
rect 21198 199448 22226 199594
rect 22394 199448 23422 199594
rect 23590 199448 24618 199594
rect 24786 199448 25814 199594
rect 25982 199448 27010 199594
rect 27178 199448 28298 199594
rect 28466 199448 29494 199594
rect 29662 199448 30690 199594
rect 30858 199448 31886 199594
rect 32054 199448 33082 199594
rect 33250 199448 34278 199594
rect 34446 199448 35474 199594
rect 35642 199448 36762 199594
rect 36930 199448 37958 199594
rect 38126 199448 39154 199594
rect 39322 199448 40350 199594
rect 40518 199448 41546 199594
rect 41714 199448 42742 199594
rect 42910 199448 43938 199594
rect 44106 199448 45134 199594
rect 45302 199448 46422 199594
rect 46590 199448 47618 199594
rect 47786 199448 48814 199594
rect 48982 199448 50010 199594
rect 50178 199448 51206 199594
rect 51374 199448 52402 199594
rect 52570 199448 53598 199594
rect 53766 199448 54886 199594
rect 55054 199448 56082 199594
rect 56250 199448 57278 199594
rect 57446 199448 58474 199594
rect 58642 199448 59670 199594
rect 59838 199448 60866 199594
rect 61034 199448 62062 199594
rect 62230 199448 63258 199594
rect 63426 199448 64546 199594
rect 64714 199448 65742 199594
rect 65910 199448 66938 199594
rect 67106 199448 68134 199594
rect 68302 199448 69330 199594
rect 69498 199448 70526 199594
rect 70694 199448 71722 199594
rect 71890 199448 73010 199594
rect 73178 199448 74206 199594
rect 74374 199448 75402 199594
rect 75570 199448 76598 199594
rect 76766 199448 77794 199594
rect 77962 199448 78990 199594
rect 79158 199448 80186 199594
rect 80354 199448 81382 199594
rect 81550 199448 82670 199594
rect 82838 199448 83866 199594
rect 84034 199448 85062 199594
rect 85230 199448 86258 199594
rect 86426 199448 87454 199594
rect 87622 199448 88650 199594
rect 88818 199448 89846 199594
rect 90014 199448 91134 199594
rect 91302 199448 92330 199594
rect 92498 199448 93526 199594
rect 93694 199448 94722 199594
rect 94890 199448 95918 199594
rect 96086 199448 97114 199594
rect 97282 199448 98310 199594
rect 98478 199448 99598 199594
rect 99766 199448 100794 199594
rect 100962 199448 101990 199594
rect 102158 199448 103186 199594
rect 103354 199448 104382 199594
rect 104550 199448 105578 199594
rect 105746 199448 106774 199594
rect 106942 199448 107970 199594
rect 108138 199448 109258 199594
rect 109426 199448 110454 199594
rect 110622 199448 111650 199594
rect 111818 199448 112846 199594
rect 113014 199448 114042 199594
rect 114210 199448 115238 199594
rect 115406 199448 116434 199594
rect 116602 199448 117722 199594
rect 117890 199448 118918 199594
rect 119086 199448 120114 199594
rect 120282 199448 121310 199594
rect 121478 199448 122506 199594
rect 122674 199448 123702 199594
rect 123870 199448 124898 199594
rect 125066 199448 126094 199594
rect 126262 199448 127382 199594
rect 127550 199448 128578 199594
rect 128746 199448 129774 199594
rect 129942 199448 130970 199594
rect 131138 199448 132166 199594
rect 132334 199448 133362 199594
rect 133530 199448 134558 199594
rect 134726 199448 135846 199594
rect 136014 199448 137042 199594
rect 137210 199448 138238 199594
rect 138406 199448 139434 199594
rect 139602 199448 140630 199594
rect 140798 199448 141826 199594
rect 141994 199448 143022 199594
rect 143190 199448 144218 199594
rect 144386 199448 145506 199594
rect 145674 199448 146702 199594
rect 146870 199448 147898 199594
rect 148066 199448 149094 199594
rect 149262 199448 150290 199594
rect 150458 199448 151486 199594
rect 151654 199448 152682 199594
rect 152850 199448 153970 199594
rect 154138 199448 155166 199594
rect 155334 199448 156362 199594
rect 156530 199448 157558 199594
rect 157726 199448 158754 199594
rect 158922 199448 159950 199594
rect 160118 199448 161146 199594
rect 161314 199448 162342 199594
rect 162510 199448 163630 199594
rect 163798 199448 164826 199594
rect 164994 199448 166022 199594
rect 166190 199448 167218 199594
rect 167386 199448 168414 199594
rect 168582 199448 169610 199594
rect 169778 199448 170806 199594
rect 170974 199448 172094 199594
rect 172262 199448 173290 199594
rect 173458 199448 174486 199594
rect 174654 199448 175682 199594
rect 175850 199448 176878 199594
rect 177046 199448 178074 199594
rect 178242 199448 179270 199594
rect 179438 199448 180466 199594
rect 180634 199448 181754 199594
rect 181922 199448 182950 199594
rect 183118 199448 184146 199594
rect 184314 199448 185342 199594
rect 185510 199448 186538 199594
rect 186706 199448 187734 199594
rect 187902 199448 188930 199594
rect 189098 199448 190218 199594
rect 190386 199448 191414 199594
rect 191582 199448 192610 199594
rect 192778 199448 193806 199594
rect 193974 199448 195002 199594
rect 195170 199448 196198 199594
rect 196366 199448 197394 199594
rect 197562 199448 197780 199594
rect 18 856 197780 199448
rect 18 614 606 856
rect 774 614 1986 856
rect 2154 614 3366 856
rect 3534 614 4746 856
rect 4914 614 6126 856
rect 6294 614 7506 856
rect 7674 614 8886 856
rect 9054 614 10266 856
rect 10434 614 11646 856
rect 11814 614 13026 856
rect 13194 614 14406 856
rect 14574 614 15786 856
rect 15954 614 17166 856
rect 17334 614 18546 856
rect 18714 614 19926 856
rect 20094 614 21306 856
rect 21474 614 22778 856
rect 22946 614 24158 856
rect 24326 614 25538 856
rect 25706 614 26918 856
rect 27086 614 28298 856
rect 28466 614 29678 856
rect 29846 614 31058 856
rect 31226 614 32438 856
rect 32606 614 33818 856
rect 33986 614 35198 856
rect 35366 614 36578 856
rect 36746 614 37958 856
rect 38126 614 39338 856
rect 39506 614 40718 856
rect 40886 614 42098 856
rect 42266 614 43478 856
rect 43646 614 44950 856
rect 45118 614 46330 856
rect 46498 614 47710 856
rect 47878 614 49090 856
rect 49258 614 50470 856
rect 50638 614 51850 856
rect 52018 614 53230 856
rect 53398 614 54610 856
rect 54778 614 55990 856
rect 56158 614 57370 856
rect 57538 614 58750 856
rect 58918 614 60130 856
rect 60298 614 61510 856
rect 61678 614 62890 856
rect 63058 614 64270 856
rect 64438 614 65650 856
rect 65818 614 67122 856
rect 67290 614 68502 856
rect 68670 614 69882 856
rect 70050 614 71262 856
rect 71430 614 72642 856
rect 72810 614 74022 856
rect 74190 614 75402 856
rect 75570 614 76782 856
rect 76950 614 78162 856
rect 78330 614 79542 856
rect 79710 614 80922 856
rect 81090 614 82302 856
rect 82470 614 83682 856
rect 83850 614 85062 856
rect 85230 614 86442 856
rect 86610 614 87822 856
rect 87990 614 89294 856
rect 89462 614 90674 856
rect 90842 614 92054 856
rect 92222 614 93434 856
rect 93602 614 94814 856
rect 94982 614 96194 856
rect 96362 614 97574 856
rect 97742 614 98954 856
rect 99122 614 100334 856
rect 100502 614 101714 856
rect 101882 614 103094 856
rect 103262 614 104474 856
rect 104642 614 105854 856
rect 106022 614 107234 856
rect 107402 614 108614 856
rect 108782 614 109994 856
rect 110162 614 111466 856
rect 111634 614 112846 856
rect 113014 614 114226 856
rect 114394 614 115606 856
rect 115774 614 116986 856
rect 117154 614 118366 856
rect 118534 614 119746 856
rect 119914 614 121126 856
rect 121294 614 122506 856
rect 122674 614 123886 856
rect 124054 614 125266 856
rect 125434 614 126646 856
rect 126814 614 128026 856
rect 128194 614 129406 856
rect 129574 614 130786 856
rect 130954 614 132166 856
rect 132334 614 133638 856
rect 133806 614 135018 856
rect 135186 614 136398 856
rect 136566 614 137778 856
rect 137946 614 139158 856
rect 139326 614 140538 856
rect 140706 614 141918 856
rect 142086 614 143298 856
rect 143466 614 144678 856
rect 144846 614 146058 856
rect 146226 614 147438 856
rect 147606 614 148818 856
rect 148986 614 150198 856
rect 150366 614 151578 856
rect 151746 614 152958 856
rect 153126 614 154338 856
rect 154506 614 155810 856
rect 155978 614 157190 856
rect 157358 614 158570 856
rect 158738 614 159950 856
rect 160118 614 161330 856
rect 161498 614 162710 856
rect 162878 614 164090 856
rect 164258 614 165470 856
rect 165638 614 166850 856
rect 167018 614 168230 856
rect 168398 614 169610 856
rect 169778 614 170990 856
rect 171158 614 172370 856
rect 172538 614 173750 856
rect 173918 614 175130 856
rect 175298 614 176510 856
rect 176678 614 177982 856
rect 178150 614 179362 856
rect 179530 614 180742 856
rect 180910 614 182122 856
rect 182290 614 183502 856
rect 183670 614 184882 856
rect 185050 614 186262 856
rect 186430 614 187642 856
rect 187810 614 189022 856
rect 189190 614 190402 856
rect 190570 614 191782 856
rect 191950 614 193162 856
rect 193330 614 194542 856
rect 194710 614 195922 856
rect 196090 614 197302 856
rect 197470 614 197780 856
<< metal3 >>
rect 0 197480 800 197600
rect 197360 197616 198160 197736
rect 197360 192448 198160 192568
rect 0 192040 800 192160
rect 197360 187280 198160 187400
rect 0 186600 800 186720
rect 197360 182112 198160 182232
rect 0 181160 800 181280
rect 197360 177080 198160 177200
rect 0 175720 800 175840
rect 197360 171912 198160 172032
rect 0 170416 800 170536
rect 197360 166744 198160 166864
rect 0 164976 800 165096
rect 197360 161576 198160 161696
rect 0 159536 800 159656
rect 197360 156544 198160 156664
rect 0 154096 800 154216
rect 197360 151376 198160 151496
rect 0 148656 800 148776
rect 197360 146208 198160 146328
rect 0 143352 800 143472
rect 197360 141040 198160 141160
rect 0 137912 800 138032
rect 197360 136008 198160 136128
rect 0 132472 800 132592
rect 197360 130840 198160 130960
rect 0 127032 800 127152
rect 197360 125672 198160 125792
rect 0 121592 800 121712
rect 197360 120504 198160 120624
rect 0 116288 800 116408
rect 197360 115336 198160 115456
rect 0 110848 800 110968
rect 197360 110304 198160 110424
rect 0 105408 800 105528
rect 197360 105136 198160 105256
rect 0 99968 800 100088
rect 197360 99968 198160 100088
rect 197360 94800 198160 94920
rect 0 94528 800 94648
rect 197360 89768 198160 89888
rect 0 89088 800 89208
rect 197360 84600 198160 84720
rect 0 83784 800 83904
rect 197360 79432 198160 79552
rect 0 78344 800 78464
rect 197360 74264 198160 74384
rect 0 72904 800 73024
rect 197360 69232 198160 69352
rect 0 67464 800 67584
rect 197360 64064 198160 64184
rect 0 62024 800 62144
rect 197360 58896 198160 59016
rect 0 56720 800 56840
rect 197360 53728 198160 53848
rect 0 51280 800 51400
rect 197360 48560 198160 48680
rect 0 45840 800 45960
rect 197360 43528 198160 43648
rect 0 40400 800 40520
rect 197360 38360 198160 38480
rect 0 34960 800 35080
rect 197360 33192 198160 33312
rect 0 29656 800 29776
rect 197360 28024 198160 28144
rect 0 24216 800 24336
rect 197360 22992 198160 23112
rect 0 18776 800 18896
rect 197360 17824 198160 17944
rect 0 13336 800 13456
rect 197360 12656 198160 12776
rect 0 7896 800 8016
rect 197360 7488 198160 7608
rect 0 2592 800 2712
rect 197360 2456 198160 2576
<< obsm3 >>
rect 13 197816 197695 198253
rect 13 197680 197280 197816
rect 880 197536 197280 197680
rect 880 197400 197695 197536
rect 13 192648 197695 197400
rect 13 192368 197280 192648
rect 13 192240 197695 192368
rect 880 191960 197695 192240
rect 13 187480 197695 191960
rect 13 187200 197280 187480
rect 13 186800 197695 187200
rect 880 186520 197695 186800
rect 13 182312 197695 186520
rect 13 182032 197280 182312
rect 13 181360 197695 182032
rect 880 181080 197695 181360
rect 13 177280 197695 181080
rect 13 177000 197280 177280
rect 13 175920 197695 177000
rect 880 175640 197695 175920
rect 13 172112 197695 175640
rect 13 171832 197280 172112
rect 13 170616 197695 171832
rect 880 170336 197695 170616
rect 13 166944 197695 170336
rect 13 166664 197280 166944
rect 13 165176 197695 166664
rect 880 164896 197695 165176
rect 13 161776 197695 164896
rect 13 161496 197280 161776
rect 13 159736 197695 161496
rect 880 159456 197695 159736
rect 13 156744 197695 159456
rect 13 156464 197280 156744
rect 13 154296 197695 156464
rect 880 154016 197695 154296
rect 13 151576 197695 154016
rect 13 151296 197280 151576
rect 13 148856 197695 151296
rect 880 148576 197695 148856
rect 13 146408 197695 148576
rect 13 146128 197280 146408
rect 13 143552 197695 146128
rect 880 143272 197695 143552
rect 13 141240 197695 143272
rect 13 140960 197280 141240
rect 13 138112 197695 140960
rect 880 137832 197695 138112
rect 13 136208 197695 137832
rect 13 135928 197280 136208
rect 13 132672 197695 135928
rect 880 132392 197695 132672
rect 13 131040 197695 132392
rect 13 130760 197280 131040
rect 13 127232 197695 130760
rect 880 126952 197695 127232
rect 13 125872 197695 126952
rect 13 125592 197280 125872
rect 13 121792 197695 125592
rect 880 121512 197695 121792
rect 13 120704 197695 121512
rect 13 120424 197280 120704
rect 13 116488 197695 120424
rect 880 116208 197695 116488
rect 13 115536 197695 116208
rect 13 115256 197280 115536
rect 13 111048 197695 115256
rect 880 110768 197695 111048
rect 13 110504 197695 110768
rect 13 110224 197280 110504
rect 13 105608 197695 110224
rect 880 105336 197695 105608
rect 880 105328 197280 105336
rect 13 105056 197280 105328
rect 13 100168 197695 105056
rect 880 99888 197280 100168
rect 13 95000 197695 99888
rect 13 94728 197280 95000
rect 880 94720 197280 94728
rect 880 94448 197695 94720
rect 13 89968 197695 94448
rect 13 89688 197280 89968
rect 13 89288 197695 89688
rect 880 89008 197695 89288
rect 13 84800 197695 89008
rect 13 84520 197280 84800
rect 13 83984 197695 84520
rect 880 83704 197695 83984
rect 13 79632 197695 83704
rect 13 79352 197280 79632
rect 13 78544 197695 79352
rect 880 78264 197695 78544
rect 13 74464 197695 78264
rect 13 74184 197280 74464
rect 13 73104 197695 74184
rect 880 72824 197695 73104
rect 13 69432 197695 72824
rect 13 69152 197280 69432
rect 13 67664 197695 69152
rect 880 67384 197695 67664
rect 13 64264 197695 67384
rect 13 63984 197280 64264
rect 13 62224 197695 63984
rect 880 61944 197695 62224
rect 13 59096 197695 61944
rect 13 58816 197280 59096
rect 13 56920 197695 58816
rect 880 56640 197695 56920
rect 13 53928 197695 56640
rect 13 53648 197280 53928
rect 13 51480 197695 53648
rect 880 51200 197695 51480
rect 13 48760 197695 51200
rect 13 48480 197280 48760
rect 13 46040 197695 48480
rect 880 45760 197695 46040
rect 13 43728 197695 45760
rect 13 43448 197280 43728
rect 13 40600 197695 43448
rect 880 40320 197695 40600
rect 13 38560 197695 40320
rect 13 38280 197280 38560
rect 13 35160 197695 38280
rect 880 34880 197695 35160
rect 13 33392 197695 34880
rect 13 33112 197280 33392
rect 13 29856 197695 33112
rect 880 29576 197695 29856
rect 13 28224 197695 29576
rect 13 27944 197280 28224
rect 13 24416 197695 27944
rect 880 24136 197695 24416
rect 13 23192 197695 24136
rect 13 22912 197280 23192
rect 13 18976 197695 22912
rect 880 18696 197695 18976
rect 13 18024 197695 18696
rect 13 17744 197280 18024
rect 13 13536 197695 17744
rect 880 13256 197695 13536
rect 13 12856 197695 13256
rect 13 12576 197280 12856
rect 13 8096 197695 12576
rect 880 7816 197695 8096
rect 13 7688 197695 7816
rect 13 7408 197280 7688
rect 13 2792 197695 7408
rect 880 2656 197695 2792
rect 880 2512 197280 2656
rect 13 2376 197280 2512
rect 13 1259 197695 2376
<< metal4 >>
rect 4208 2128 4528 198064
rect 19568 2128 19888 198064
rect 34928 2128 35248 198064
rect 50288 2128 50608 198064
rect 65648 2128 65968 198064
rect 81008 2128 81328 198064
rect 96368 2128 96688 198064
rect 111728 2128 112048 198064
rect 127088 2128 127408 198064
rect 142448 2128 142768 198064
rect 157808 2128 158128 198064
rect 173168 2128 173488 198064
rect 188528 2128 188848 198064
<< obsm4 >>
rect 23979 198144 192589 198253
rect 23979 2048 34848 198144
rect 35328 2048 50208 198144
rect 50688 2048 65568 198144
rect 66048 2048 80928 198144
rect 81408 2048 96288 198144
rect 96768 2048 111648 198144
rect 112128 2048 127008 198144
rect 127488 2048 142368 198144
rect 142848 2048 157728 198144
rect 158208 2048 173088 198144
rect 173568 2048 188448 198144
rect 188928 2048 192589 198144
rect 23979 1259 192589 2048
<< labels >>
rlabel metal3 s 197360 2456 198160 2576 6 clk_i
port 1 nsew signal input
rlabel metal3 s 197360 7488 198160 7608 6 i_dout0[0]
port 2 nsew signal input
rlabel metal3 s 197360 94800 198160 94920 6 i_dout0[10]
port 3 nsew signal input
rlabel metal3 s 197360 99968 198160 100088 6 i_dout0[11]
port 4 nsew signal input
rlabel metal3 s 197360 110304 198160 110424 6 i_dout0[12]
port 5 nsew signal input
rlabel metal3 s 0 83784 800 83904 6 i_dout0[13]
port 6 nsew signal input
rlabel metal2 s 170862 199504 170918 200304 6 i_dout0[14]
port 7 nsew signal input
rlabel metal2 s 173346 199504 173402 200304 6 i_dout0[15]
port 8 nsew signal input
rlabel metal3 s 0 105408 800 105528 6 i_dout0[16]
port 9 nsew signal input
rlabel metal2 s 176934 199504 176990 200304 6 i_dout0[17]
port 10 nsew signal input
rlabel metal3 s 197360 130840 198160 130960 6 i_dout0[18]
port 11 nsew signal input
rlabel metal3 s 0 121592 800 121712 6 i_dout0[19]
port 12 nsew signal input
rlabel metal2 s 153014 0 153070 800 6 i_dout0[1]
port 13 nsew signal input
rlabel metal3 s 197360 141040 198160 141160 6 i_dout0[20]
port 14 nsew signal input
rlabel metal2 s 184202 199504 184258 200304 6 i_dout0[21]
port 15 nsew signal input
rlabel metal2 s 185398 199504 185454 200304 6 i_dout0[22]
port 16 nsew signal input
rlabel metal3 s 0 143352 800 143472 6 i_dout0[23]
port 17 nsew signal input
rlabel metal2 s 186594 199504 186650 200304 6 i_dout0[24]
port 18 nsew signal input
rlabel metal2 s 187790 199504 187846 200304 6 i_dout0[25]
port 19 nsew signal input
rlabel metal2 s 191470 199504 191526 200304 6 i_dout0[26]
port 20 nsew signal input
rlabel metal2 s 191838 0 191894 800 6 i_dout0[27]
port 21 nsew signal input
rlabel metal3 s 197360 187280 198160 187400 6 i_dout0[28]
port 22 nsew signal input
rlabel metal2 s 194598 0 194654 800 6 i_dout0[29]
port 23 nsew signal input
rlabel metal2 s 160006 0 160062 800 6 i_dout0[2]
port 24 nsew signal input
rlabel metal3 s 0 192040 800 192160 6 i_dout0[30]
port 25 nsew signal input
rlabel metal3 s 0 197480 800 197600 6 i_dout0[31]
port 26 nsew signal input
rlabel metal3 s 0 24216 800 24336 6 i_dout0[3]
port 27 nsew signal input
rlabel metal3 s 197360 53728 198160 53848 6 i_dout0[4]
port 28 nsew signal input
rlabel metal2 s 150346 199504 150402 200304 6 i_dout0[5]
port 29 nsew signal input
rlabel metal3 s 197360 74264 198160 74384 6 i_dout0[6]
port 30 nsew signal input
rlabel metal2 s 158810 199504 158866 200304 6 i_dout0[7]
port 31 nsew signal input
rlabel metal2 s 173806 0 173862 800 6 i_dout0[8]
port 32 nsew signal input
rlabel metal2 s 176566 0 176622 800 6 i_dout0[9]
port 33 nsew signal input
rlabel metal2 s 141882 199504 141938 200304 6 i_dout0_1[0]
port 34 nsew signal input
rlabel metal3 s 197360 89768 198160 89888 6 i_dout0_1[10]
port 35 nsew signal input
rlabel metal2 s 179418 0 179474 800 6 i_dout0_1[11]
port 36 nsew signal input
rlabel metal2 s 166078 199504 166134 200304 6 i_dout0_1[12]
port 37 nsew signal input
rlabel metal3 s 0 78344 800 78464 6 i_dout0_1[13]
port 38 nsew signal input
rlabel metal3 s 197360 120504 198160 120624 6 i_dout0_1[14]
port 39 nsew signal input
rlabel metal2 s 182178 0 182234 800 6 i_dout0_1[15]
port 40 nsew signal input
rlabel metal2 s 174542 199504 174598 200304 6 i_dout0_1[16]
port 41 nsew signal input
rlabel metal2 s 175738 199504 175794 200304 6 i_dout0_1[17]
port 42 nsew signal input
rlabel metal2 s 180522 199504 180578 200304 6 i_dout0_1[18]
port 43 nsew signal input
rlabel metal2 s 183006 199504 183062 200304 6 i_dout0_1[19]
port 44 nsew signal input
rlabel metal3 s 0 13336 800 13456 6 i_dout0_1[1]
port 45 nsew signal input
rlabel metal2 s 183558 0 183614 800 6 i_dout0_1[20]
port 46 nsew signal input
rlabel metal3 s 197360 146208 198160 146328 6 i_dout0_1[21]
port 47 nsew signal input
rlabel metal3 s 197360 151376 198160 151496 6 i_dout0_1[22]
port 48 nsew signal input
rlabel metal2 s 189078 0 189134 800 6 i_dout0_1[23]
port 49 nsew signal input
rlabel metal3 s 197360 166744 198160 166864 6 i_dout0_1[24]
port 50 nsew signal input
rlabel metal2 s 190458 0 190514 800 6 i_dout0_1[25]
port 51 nsew signal input
rlabel metal2 s 190274 199504 190330 200304 6 i_dout0_1[26]
port 52 nsew signal input
rlabel metal3 s 197360 182112 198160 182232 6 i_dout0_1[27]
port 53 nsew signal input
rlabel metal2 s 193862 199504 193918 200304 6 i_dout0_1[28]
port 54 nsew signal input
rlabel metal3 s 0 181160 800 181280 6 i_dout0_1[29]
port 55 nsew signal input
rlabel metal2 s 158626 0 158682 800 6 i_dout0_1[2]
port 56 nsew signal input
rlabel metal2 s 196254 199504 196310 200304 6 i_dout0_1[30]
port 57 nsew signal input
rlabel metal2 s 197358 0 197414 800 6 i_dout0_1[31]
port 58 nsew signal input
rlabel metal3 s 197360 38360 198160 38480 6 i_dout0_1[3]
port 59 nsew signal input
rlabel metal2 s 149150 199504 149206 200304 6 i_dout0_1[4]
port 60 nsew signal input
rlabel metal3 s 197360 69232 198160 69352 6 i_dout0_1[5]
port 61 nsew signal input
rlabel metal2 s 154026 199504 154082 200304 6 i_dout0_1[6]
port 62 nsew signal input
rlabel metal2 s 157614 199504 157670 200304 6 i_dout0_1[7]
port 63 nsew signal input
rlabel metal2 s 161202 199504 161258 200304 6 i_dout0_1[8]
port 64 nsew signal input
rlabel metal2 s 163686 199504 163742 200304 6 i_dout0_1[9]
port 65 nsew signal input
rlabel metal2 s 570 199504 626 200304 6 io_in[0]
port 66 nsew signal input
rlabel metal2 s 36818 199504 36874 200304 6 io_in[10]
port 67 nsew signal input
rlabel metal2 s 40406 199504 40462 200304 6 io_in[11]
port 68 nsew signal input
rlabel metal2 s 43994 199504 44050 200304 6 io_in[12]
port 69 nsew signal input
rlabel metal2 s 47674 199504 47730 200304 6 io_in[13]
port 70 nsew signal input
rlabel metal2 s 51262 199504 51318 200304 6 io_in[14]
port 71 nsew signal input
rlabel metal2 s 54942 199504 54998 200304 6 io_in[15]
port 72 nsew signal input
rlabel metal2 s 58530 199504 58586 200304 6 io_in[16]
port 73 nsew signal input
rlabel metal2 s 62118 199504 62174 200304 6 io_in[17]
port 74 nsew signal input
rlabel metal2 s 65798 199504 65854 200304 6 io_in[18]
port 75 nsew signal input
rlabel metal2 s 69386 199504 69442 200304 6 io_in[19]
port 76 nsew signal input
rlabel metal2 s 4158 199504 4214 200304 6 io_in[1]
port 77 nsew signal input
rlabel metal2 s 73066 199504 73122 200304 6 io_in[20]
port 78 nsew signal input
rlabel metal2 s 76654 199504 76710 200304 6 io_in[21]
port 79 nsew signal input
rlabel metal2 s 80242 199504 80298 200304 6 io_in[22]
port 80 nsew signal input
rlabel metal2 s 83922 199504 83978 200304 6 io_in[23]
port 81 nsew signal input
rlabel metal2 s 87510 199504 87566 200304 6 io_in[24]
port 82 nsew signal input
rlabel metal2 s 91190 199504 91246 200304 6 io_in[25]
port 83 nsew signal input
rlabel metal2 s 94778 199504 94834 200304 6 io_in[26]
port 84 nsew signal input
rlabel metal2 s 98366 199504 98422 200304 6 io_in[27]
port 85 nsew signal input
rlabel metal2 s 102046 199504 102102 200304 6 io_in[28]
port 86 nsew signal input
rlabel metal2 s 105634 199504 105690 200304 6 io_in[29]
port 87 nsew signal input
rlabel metal2 s 7746 199504 7802 200304 6 io_in[2]
port 88 nsew signal input
rlabel metal2 s 109314 199504 109370 200304 6 io_in[30]
port 89 nsew signal input
rlabel metal2 s 112902 199504 112958 200304 6 io_in[31]
port 90 nsew signal input
rlabel metal2 s 116490 199504 116546 200304 6 io_in[32]
port 91 nsew signal input
rlabel metal2 s 120170 199504 120226 200304 6 io_in[33]
port 92 nsew signal input
rlabel metal2 s 123758 199504 123814 200304 6 io_in[34]
port 93 nsew signal input
rlabel metal2 s 127438 199504 127494 200304 6 io_in[35]
port 94 nsew signal input
rlabel metal2 s 131026 199504 131082 200304 6 io_in[36]
port 95 nsew signal input
rlabel metal2 s 134614 199504 134670 200304 6 io_in[37]
port 96 nsew signal input
rlabel metal2 s 11426 199504 11482 200304 6 io_in[3]
port 97 nsew signal input
rlabel metal2 s 15014 199504 15070 200304 6 io_in[4]
port 98 nsew signal input
rlabel metal2 s 18694 199504 18750 200304 6 io_in[5]
port 99 nsew signal input
rlabel metal2 s 22282 199504 22338 200304 6 io_in[6]
port 100 nsew signal input
rlabel metal2 s 25870 199504 25926 200304 6 io_in[7]
port 101 nsew signal input
rlabel metal2 s 29550 199504 29606 200304 6 io_in[8]
port 102 nsew signal input
rlabel metal2 s 33138 199504 33194 200304 6 io_in[9]
port 103 nsew signal input
rlabel metal2 s 1766 199504 1822 200304 6 io_oeb[0]
port 104 nsew signal output
rlabel metal2 s 38014 199504 38070 200304 6 io_oeb[10]
port 105 nsew signal output
rlabel metal2 s 41602 199504 41658 200304 6 io_oeb[11]
port 106 nsew signal output
rlabel metal2 s 45190 199504 45246 200304 6 io_oeb[12]
port 107 nsew signal output
rlabel metal2 s 48870 199504 48926 200304 6 io_oeb[13]
port 108 nsew signal output
rlabel metal2 s 52458 199504 52514 200304 6 io_oeb[14]
port 109 nsew signal output
rlabel metal2 s 56138 199504 56194 200304 6 io_oeb[15]
port 110 nsew signal output
rlabel metal2 s 59726 199504 59782 200304 6 io_oeb[16]
port 111 nsew signal output
rlabel metal2 s 63314 199504 63370 200304 6 io_oeb[17]
port 112 nsew signal output
rlabel metal2 s 66994 199504 67050 200304 6 io_oeb[18]
port 113 nsew signal output
rlabel metal2 s 70582 199504 70638 200304 6 io_oeb[19]
port 114 nsew signal output
rlabel metal2 s 5354 199504 5410 200304 6 io_oeb[1]
port 115 nsew signal output
rlabel metal2 s 74262 199504 74318 200304 6 io_oeb[20]
port 116 nsew signal output
rlabel metal2 s 77850 199504 77906 200304 6 io_oeb[21]
port 117 nsew signal output
rlabel metal2 s 81438 199504 81494 200304 6 io_oeb[22]
port 118 nsew signal output
rlabel metal2 s 85118 199504 85174 200304 6 io_oeb[23]
port 119 nsew signal output
rlabel metal2 s 88706 199504 88762 200304 6 io_oeb[24]
port 120 nsew signal output
rlabel metal2 s 92386 199504 92442 200304 6 io_oeb[25]
port 121 nsew signal output
rlabel metal2 s 95974 199504 96030 200304 6 io_oeb[26]
port 122 nsew signal output
rlabel metal2 s 99654 199504 99710 200304 6 io_oeb[27]
port 123 nsew signal output
rlabel metal2 s 103242 199504 103298 200304 6 io_oeb[28]
port 124 nsew signal output
rlabel metal2 s 106830 199504 106886 200304 6 io_oeb[29]
port 125 nsew signal output
rlabel metal2 s 8942 199504 8998 200304 6 io_oeb[2]
port 126 nsew signal output
rlabel metal2 s 110510 199504 110566 200304 6 io_oeb[30]
port 127 nsew signal output
rlabel metal2 s 114098 199504 114154 200304 6 io_oeb[31]
port 128 nsew signal output
rlabel metal2 s 117778 199504 117834 200304 6 io_oeb[32]
port 129 nsew signal output
rlabel metal2 s 121366 199504 121422 200304 6 io_oeb[33]
port 130 nsew signal output
rlabel metal2 s 124954 199504 125010 200304 6 io_oeb[34]
port 131 nsew signal output
rlabel metal2 s 128634 199504 128690 200304 6 io_oeb[35]
port 132 nsew signal output
rlabel metal2 s 132222 199504 132278 200304 6 io_oeb[36]
port 133 nsew signal output
rlabel metal2 s 135902 199504 135958 200304 6 io_oeb[37]
port 134 nsew signal output
rlabel metal2 s 12622 199504 12678 200304 6 io_oeb[3]
port 135 nsew signal output
rlabel metal2 s 16210 199504 16266 200304 6 io_oeb[4]
port 136 nsew signal output
rlabel metal2 s 19890 199504 19946 200304 6 io_oeb[5]
port 137 nsew signal output
rlabel metal2 s 23478 199504 23534 200304 6 io_oeb[6]
port 138 nsew signal output
rlabel metal2 s 27066 199504 27122 200304 6 io_oeb[7]
port 139 nsew signal output
rlabel metal2 s 30746 199504 30802 200304 6 io_oeb[8]
port 140 nsew signal output
rlabel metal2 s 34334 199504 34390 200304 6 io_oeb[9]
port 141 nsew signal output
rlabel metal2 s 2962 199504 3018 200304 6 io_out[0]
port 142 nsew signal output
rlabel metal2 s 39210 199504 39266 200304 6 io_out[10]
port 143 nsew signal output
rlabel metal2 s 42798 199504 42854 200304 6 io_out[11]
port 144 nsew signal output
rlabel metal2 s 46478 199504 46534 200304 6 io_out[12]
port 145 nsew signal output
rlabel metal2 s 50066 199504 50122 200304 6 io_out[13]
port 146 nsew signal output
rlabel metal2 s 53654 199504 53710 200304 6 io_out[14]
port 147 nsew signal output
rlabel metal2 s 57334 199504 57390 200304 6 io_out[15]
port 148 nsew signal output
rlabel metal2 s 60922 199504 60978 200304 6 io_out[16]
port 149 nsew signal output
rlabel metal2 s 64602 199504 64658 200304 6 io_out[17]
port 150 nsew signal output
rlabel metal2 s 68190 199504 68246 200304 6 io_out[18]
port 151 nsew signal output
rlabel metal2 s 71778 199504 71834 200304 6 io_out[19]
port 152 nsew signal output
rlabel metal2 s 6550 199504 6606 200304 6 io_out[1]
port 153 nsew signal output
rlabel metal2 s 75458 199504 75514 200304 6 io_out[20]
port 154 nsew signal output
rlabel metal2 s 79046 199504 79102 200304 6 io_out[21]
port 155 nsew signal output
rlabel metal2 s 82726 199504 82782 200304 6 io_out[22]
port 156 nsew signal output
rlabel metal2 s 86314 199504 86370 200304 6 io_out[23]
port 157 nsew signal output
rlabel metal2 s 89902 199504 89958 200304 6 io_out[24]
port 158 nsew signal output
rlabel metal2 s 93582 199504 93638 200304 6 io_out[25]
port 159 nsew signal output
rlabel metal2 s 97170 199504 97226 200304 6 io_out[26]
port 160 nsew signal output
rlabel metal2 s 100850 199504 100906 200304 6 io_out[27]
port 161 nsew signal output
rlabel metal2 s 104438 199504 104494 200304 6 io_out[28]
port 162 nsew signal output
rlabel metal2 s 108026 199504 108082 200304 6 io_out[29]
port 163 nsew signal output
rlabel metal2 s 10230 199504 10286 200304 6 io_out[2]
port 164 nsew signal output
rlabel metal2 s 111706 199504 111762 200304 6 io_out[30]
port 165 nsew signal output
rlabel metal2 s 115294 199504 115350 200304 6 io_out[31]
port 166 nsew signal output
rlabel metal2 s 118974 199504 119030 200304 6 io_out[32]
port 167 nsew signal output
rlabel metal2 s 122562 199504 122618 200304 6 io_out[33]
port 168 nsew signal output
rlabel metal2 s 126150 199504 126206 200304 6 io_out[34]
port 169 nsew signal output
rlabel metal2 s 129830 199504 129886 200304 6 io_out[35]
port 170 nsew signal output
rlabel metal2 s 133418 199504 133474 200304 6 io_out[36]
port 171 nsew signal output
rlabel metal2 s 137098 199504 137154 200304 6 io_out[37]
port 172 nsew signal output
rlabel metal2 s 13818 199504 13874 200304 6 io_out[3]
port 173 nsew signal output
rlabel metal2 s 17406 199504 17462 200304 6 io_out[4]
port 174 nsew signal output
rlabel metal2 s 21086 199504 21142 200304 6 io_out[5]
port 175 nsew signal output
rlabel metal2 s 24674 199504 24730 200304 6 io_out[6]
port 176 nsew signal output
rlabel metal2 s 28354 199504 28410 200304 6 io_out[7]
port 177 nsew signal output
rlabel metal2 s 31942 199504 31998 200304 6 io_out[8]
port 178 nsew signal output
rlabel metal2 s 35530 199504 35586 200304 6 io_out[9]
port 179 nsew signal output
rlabel metal2 s 147494 0 147550 800 6 irq[0]
port 180 nsew signal output
rlabel metal2 s 148874 0 148930 800 6 irq[1]
port 181 nsew signal output
rlabel metal2 s 150254 0 150310 800 6 irq[2]
port 182 nsew signal output
rlabel metal3 s 0 2592 800 2712 6 o_csb0
port 183 nsew signal output
rlabel metal2 s 138294 199504 138350 200304 6 o_csb0_1
port 184 nsew signal output
rlabel metal3 s 197360 12656 198160 12776 6 o_din0[0]
port 185 nsew signal output
rlabel metal2 s 164882 199504 164938 200304 6 o_din0[10]
port 186 nsew signal output
rlabel metal2 s 180798 0 180854 800 6 o_din0[11]
port 187 nsew signal output
rlabel metal2 s 167274 199504 167330 200304 6 o_din0[12]
port 188 nsew signal output
rlabel metal2 s 169666 199504 169722 200304 6 o_din0[13]
port 189 nsew signal output
rlabel metal2 s 172150 199504 172206 200304 6 o_din0[14]
port 190 nsew signal output
rlabel metal3 s 0 99968 800 100088 6 o_din0[15]
port 191 nsew signal output
rlabel metal3 s 0 110848 800 110968 6 o_din0[16]
port 192 nsew signal output
rlabel metal2 s 179326 199504 179382 200304 6 o_din0[17]
port 193 nsew signal output
rlabel metal3 s 0 116288 800 116408 6 o_din0[18]
port 194 nsew signal output
rlabel metal3 s 0 127032 800 127152 6 o_din0[19]
port 195 nsew signal output
rlabel metal2 s 155866 0 155922 800 6 o_din0[1]
port 196 nsew signal output
rlabel metal3 s 0 132472 800 132592 6 o_din0[20]
port 197 nsew signal output
rlabel metal2 s 186318 0 186374 800 6 o_din0[21]
port 198 nsew signal output
rlabel metal3 s 197360 156544 198160 156664 6 o_din0[22]
port 199 nsew signal output
rlabel metal3 s 197360 161576 198160 161696 6 o_din0[23]
port 200 nsew signal output
rlabel metal3 s 0 154096 800 154216 6 o_din0[24]
port 201 nsew signal output
rlabel metal3 s 0 159536 800 159656 6 o_din0[25]
port 202 nsew signal output
rlabel metal2 s 192666 199504 192722 200304 6 o_din0[26]
port 203 nsew signal output
rlabel metal2 s 193218 0 193274 800 6 o_din0[27]
port 204 nsew signal output
rlabel metal3 s 0 175720 800 175840 6 o_din0[28]
port 205 nsew signal output
rlabel metal2 s 195058 199504 195114 200304 6 o_din0[29]
port 206 nsew signal output
rlabel metal2 s 161386 0 161442 800 6 o_din0[2]
port 207 nsew signal output
rlabel metal3 s 197360 192448 198160 192568 6 o_din0[30]
port 208 nsew signal output
rlabel metal2 s 197450 199504 197506 200304 6 o_din0[31]
port 209 nsew signal output
rlabel metal2 s 146758 199504 146814 200304 6 o_din0[3]
port 210 nsew signal output
rlabel metal3 s 0 40400 800 40520 6 o_din0[4]
port 211 nsew signal output
rlabel metal2 s 151542 199504 151598 200304 6 o_din0[5]
port 212 nsew signal output
rlabel metal2 s 155222 199504 155278 200304 6 o_din0[6]
port 213 nsew signal output
rlabel metal2 s 172426 0 172482 800 6 o_din0[7]
port 214 nsew signal output
rlabel metal2 s 175186 0 175242 800 6 o_din0[8]
port 215 nsew signal output
rlabel metal2 s 178038 0 178094 800 6 o_din0[9]
port 216 nsew signal output
rlabel metal3 s 0 7896 800 8016 6 o_din0_1[0]
port 217 nsew signal output
rlabel metal3 s 0 72904 800 73024 6 o_din0_1[10]
port 218 nsew signal output
rlabel metal3 s 197360 105136 198160 105256 6 o_din0_1[11]
port 219 nsew signal output
rlabel metal3 s 197360 115336 198160 115456 6 o_din0_1[12]
port 220 nsew signal output
rlabel metal2 s 168470 199504 168526 200304 6 o_din0_1[13]
port 221 nsew signal output
rlabel metal3 s 0 89088 800 89208 6 o_din0_1[14]
port 222 nsew signal output
rlabel metal3 s 0 94528 800 94648 6 o_din0_1[15]
port 223 nsew signal output
rlabel metal3 s 197360 125672 198160 125792 6 o_din0_1[16]
port 224 nsew signal output
rlabel metal2 s 178130 199504 178186 200304 6 o_din0_1[17]
port 225 nsew signal output
rlabel metal2 s 181810 199504 181866 200304 6 o_din0_1[18]
port 226 nsew signal output
rlabel metal3 s 197360 136008 198160 136128 6 o_din0_1[19]
port 227 nsew signal output
rlabel metal2 s 154394 0 154450 800 6 o_din0_1[1]
port 228 nsew signal output
rlabel metal2 s 184938 0 184994 800 6 o_din0_1[20]
port 229 nsew signal output
rlabel metal3 s 0 137912 800 138032 6 o_din0_1[21]
port 230 nsew signal output
rlabel metal2 s 187698 0 187754 800 6 o_din0_1[22]
port 231 nsew signal output
rlabel metal3 s 0 148656 800 148776 6 o_din0_1[23]
port 232 nsew signal output
rlabel metal3 s 197360 171912 198160 172032 6 o_din0_1[24]
port 233 nsew signal output
rlabel metal2 s 188986 199504 189042 200304 6 o_din0_1[25]
port 234 nsew signal output
rlabel metal3 s 197360 177080 198160 177200 6 o_din0_1[26]
port 235 nsew signal output
rlabel metal3 s 0 164976 800 165096 6 o_din0_1[27]
port 236 nsew signal output
rlabel metal3 s 0 170416 800 170536 6 o_din0_1[28]
port 237 nsew signal output
rlabel metal3 s 0 186600 800 186720 6 o_din0_1[29]
port 238 nsew signal output
rlabel metal2 s 145562 199504 145618 200304 6 o_din0_1[2]
port 239 nsew signal output
rlabel metal2 s 195978 0 196034 800 6 o_din0_1[30]
port 240 nsew signal output
rlabel metal3 s 197360 197616 198160 197736 6 o_din0_1[31]
port 241 nsew signal output
rlabel metal3 s 197360 43528 198160 43648 6 o_din0_1[3]
port 242 nsew signal output
rlabel metal3 s 197360 58896 198160 59016 6 o_din0_1[4]
port 243 nsew signal output
rlabel metal3 s 0 45840 800 45960 6 o_din0_1[5]
port 244 nsew signal output
rlabel metal2 s 171046 0 171102 800 6 o_din0_1[6]
port 245 nsew signal output
rlabel metal3 s 0 51280 800 51400 6 o_din0_1[7]
port 246 nsew signal output
rlabel metal3 s 0 62024 800 62144 6 o_din0_1[8]
port 247 nsew signal output
rlabel metal3 s 0 67464 800 67584 6 o_din0_1[9]
port 248 nsew signal output
rlabel metal3 s 197360 17824 198160 17944 6 o_waddr0[0]
port 249 nsew signal output
rlabel metal2 s 157246 0 157302 800 6 o_waddr0[1]
port 250 nsew signal output
rlabel metal2 s 164146 0 164202 800 6 o_waddr0[2]
port 251 nsew signal output
rlabel metal3 s 0 29656 800 29776 6 o_waddr0[3]
port 252 nsew signal output
rlabel metal3 s 197360 64064 198160 64184 6 o_waddr0[4]
port 253 nsew signal output
rlabel metal2 s 169666 0 169722 800 6 o_waddr0[5]
port 254 nsew signal output
rlabel metal2 s 156418 199504 156474 200304 6 o_waddr0[6]
port 255 nsew signal output
rlabel metal3 s 0 56720 800 56840 6 o_waddr0[7]
port 256 nsew signal output
rlabel metal3 s 197360 84600 198160 84720 6 o_waddr0[8]
port 257 nsew signal output
rlabel metal2 s 143078 199504 143134 200304 6 o_waddr0_1[0]
port 258 nsew signal output
rlabel metal3 s 0 18776 800 18896 6 o_waddr0_1[1]
port 259 nsew signal output
rlabel metal2 s 162766 0 162822 800 6 o_waddr0_1[2]
port 260 nsew signal output
rlabel metal2 s 147954 199504 148010 200304 6 o_waddr0_1[3]
port 261 nsew signal output
rlabel metal2 s 168286 0 168342 800 6 o_waddr0_1[4]
port 262 nsew signal output
rlabel metal2 s 152738 199504 152794 200304 6 o_waddr0_1[5]
port 263 nsew signal output
rlabel metal3 s 197360 79432 198160 79552 6 o_waddr0_1[6]
port 264 nsew signal output
rlabel metal2 s 160006 199504 160062 200304 6 o_waddr0_1[7]
port 265 nsew signal output
rlabel metal2 s 162398 199504 162454 200304 6 o_waddr0_1[8]
port 266 nsew signal output
rlabel metal2 s 139490 199504 139546 200304 6 o_web0
port 267 nsew signal output
rlabel metal2 s 140686 199504 140742 200304 6 o_web0_1
port 268 nsew signal output
rlabel metal3 s 197360 22992 198160 23112 6 o_wmask0[0]
port 269 nsew signal output
rlabel metal3 s 197360 33192 198160 33312 6 o_wmask0[1]
port 270 nsew signal output
rlabel metal2 s 166906 0 166962 800 6 o_wmask0[2]
port 271 nsew signal output
rlabel metal3 s 197360 48560 198160 48680 6 o_wmask0[3]
port 272 nsew signal output
rlabel metal3 s 197360 28024 198160 28144 6 o_wmask0_1[0]
port 273 nsew signal output
rlabel metal2 s 144274 199504 144330 200304 6 o_wmask0_1[1]
port 274 nsew signal output
rlabel metal2 s 165526 0 165582 800 6 o_wmask0_1[2]
port 275 nsew signal output
rlabel metal3 s 0 34960 800 35080 6 o_wmask0_1[3]
port 276 nsew signal output
rlabel metal2 s 151634 0 151690 800 6 rst_i
port 277 nsew signal input
rlabel metal4 s 4208 2128 4528 198064 6 vccd1
port 278 nsew power input
rlabel metal4 s 34928 2128 35248 198064 6 vccd1
port 278 nsew power input
rlabel metal4 s 65648 2128 65968 198064 6 vccd1
port 278 nsew power input
rlabel metal4 s 96368 2128 96688 198064 6 vccd1
port 278 nsew power input
rlabel metal4 s 127088 2128 127408 198064 6 vccd1
port 278 nsew power input
rlabel metal4 s 157808 2128 158128 198064 6 vccd1
port 278 nsew power input
rlabel metal4 s 188528 2128 188848 198064 6 vccd1
port 278 nsew power input
rlabel metal4 s 19568 2128 19888 198064 6 vssd1
port 279 nsew ground input
rlabel metal4 s 50288 2128 50608 198064 6 vssd1
port 279 nsew ground input
rlabel metal4 s 81008 2128 81328 198064 6 vssd1
port 279 nsew ground input
rlabel metal4 s 111728 2128 112048 198064 6 vssd1
port 279 nsew ground input
rlabel metal4 s 142448 2128 142768 198064 6 vssd1
port 279 nsew ground input
rlabel metal4 s 173168 2128 173488 198064 6 vssd1
port 279 nsew ground input
rlabel metal2 s 662 0 718 800 6 wb_clk_i
port 280 nsew signal input
rlabel metal2 s 2042 0 2098 800 6 wb_rst_i
port 281 nsew signal input
rlabel metal2 s 3422 0 3478 800 6 wbs_ack_o
port 282 nsew signal output
rlabel metal2 s 8942 0 8998 800 6 wbs_adr_i[0]
port 283 nsew signal input
rlabel metal2 s 56046 0 56102 800 6 wbs_adr_i[10]
port 284 nsew signal input
rlabel metal2 s 60186 0 60242 800 6 wbs_adr_i[11]
port 285 nsew signal input
rlabel metal2 s 64326 0 64382 800 6 wbs_adr_i[12]
port 286 nsew signal input
rlabel metal2 s 68558 0 68614 800 6 wbs_adr_i[13]
port 287 nsew signal input
rlabel metal2 s 72698 0 72754 800 6 wbs_adr_i[14]
port 288 nsew signal input
rlabel metal2 s 76838 0 76894 800 6 wbs_adr_i[15]
port 289 nsew signal input
rlabel metal2 s 80978 0 81034 800 6 wbs_adr_i[16]
port 290 nsew signal input
rlabel metal2 s 85118 0 85174 800 6 wbs_adr_i[17]
port 291 nsew signal input
rlabel metal2 s 89350 0 89406 800 6 wbs_adr_i[18]
port 292 nsew signal input
rlabel metal2 s 93490 0 93546 800 6 wbs_adr_i[19]
port 293 nsew signal input
rlabel metal2 s 14462 0 14518 800 6 wbs_adr_i[1]
port 294 nsew signal input
rlabel metal2 s 97630 0 97686 800 6 wbs_adr_i[20]
port 295 nsew signal input
rlabel metal2 s 101770 0 101826 800 6 wbs_adr_i[21]
port 296 nsew signal input
rlabel metal2 s 105910 0 105966 800 6 wbs_adr_i[22]
port 297 nsew signal input
rlabel metal2 s 110050 0 110106 800 6 wbs_adr_i[23]
port 298 nsew signal input
rlabel metal2 s 114282 0 114338 800 6 wbs_adr_i[24]
port 299 nsew signal input
rlabel metal2 s 118422 0 118478 800 6 wbs_adr_i[25]
port 300 nsew signal input
rlabel metal2 s 122562 0 122618 800 6 wbs_adr_i[26]
port 301 nsew signal input
rlabel metal2 s 126702 0 126758 800 6 wbs_adr_i[27]
port 302 nsew signal input
rlabel metal2 s 130842 0 130898 800 6 wbs_adr_i[28]
port 303 nsew signal input
rlabel metal2 s 135074 0 135130 800 6 wbs_adr_i[29]
port 304 nsew signal input
rlabel metal2 s 19982 0 20038 800 6 wbs_adr_i[2]
port 305 nsew signal input
rlabel metal2 s 139214 0 139270 800 6 wbs_adr_i[30]
port 306 nsew signal input
rlabel metal2 s 143354 0 143410 800 6 wbs_adr_i[31]
port 307 nsew signal input
rlabel metal2 s 25594 0 25650 800 6 wbs_adr_i[3]
port 308 nsew signal input
rlabel metal2 s 31114 0 31170 800 6 wbs_adr_i[4]
port 309 nsew signal input
rlabel metal2 s 35254 0 35310 800 6 wbs_adr_i[5]
port 310 nsew signal input
rlabel metal2 s 39394 0 39450 800 6 wbs_adr_i[6]
port 311 nsew signal input
rlabel metal2 s 43534 0 43590 800 6 wbs_adr_i[7]
port 312 nsew signal input
rlabel metal2 s 47766 0 47822 800 6 wbs_adr_i[8]
port 313 nsew signal input
rlabel metal2 s 51906 0 51962 800 6 wbs_adr_i[9]
port 314 nsew signal input
rlabel metal2 s 4802 0 4858 800 6 wbs_cyc_i
port 315 nsew signal input
rlabel metal2 s 10322 0 10378 800 6 wbs_dat_i[0]
port 316 nsew signal input
rlabel metal2 s 57426 0 57482 800 6 wbs_dat_i[10]
port 317 nsew signal input
rlabel metal2 s 61566 0 61622 800 6 wbs_dat_i[11]
port 318 nsew signal input
rlabel metal2 s 65706 0 65762 800 6 wbs_dat_i[12]
port 319 nsew signal input
rlabel metal2 s 69938 0 69994 800 6 wbs_dat_i[13]
port 320 nsew signal input
rlabel metal2 s 74078 0 74134 800 6 wbs_dat_i[14]
port 321 nsew signal input
rlabel metal2 s 78218 0 78274 800 6 wbs_dat_i[15]
port 322 nsew signal input
rlabel metal2 s 82358 0 82414 800 6 wbs_dat_i[16]
port 323 nsew signal input
rlabel metal2 s 86498 0 86554 800 6 wbs_dat_i[17]
port 324 nsew signal input
rlabel metal2 s 90730 0 90786 800 6 wbs_dat_i[18]
port 325 nsew signal input
rlabel metal2 s 94870 0 94926 800 6 wbs_dat_i[19]
port 326 nsew signal input
rlabel metal2 s 15842 0 15898 800 6 wbs_dat_i[1]
port 327 nsew signal input
rlabel metal2 s 99010 0 99066 800 6 wbs_dat_i[20]
port 328 nsew signal input
rlabel metal2 s 103150 0 103206 800 6 wbs_dat_i[21]
port 329 nsew signal input
rlabel metal2 s 107290 0 107346 800 6 wbs_dat_i[22]
port 330 nsew signal input
rlabel metal2 s 111522 0 111578 800 6 wbs_dat_i[23]
port 331 nsew signal input
rlabel metal2 s 115662 0 115718 800 6 wbs_dat_i[24]
port 332 nsew signal input
rlabel metal2 s 119802 0 119858 800 6 wbs_dat_i[25]
port 333 nsew signal input
rlabel metal2 s 123942 0 123998 800 6 wbs_dat_i[26]
port 334 nsew signal input
rlabel metal2 s 128082 0 128138 800 6 wbs_dat_i[27]
port 335 nsew signal input
rlabel metal2 s 132222 0 132278 800 6 wbs_dat_i[28]
port 336 nsew signal input
rlabel metal2 s 136454 0 136510 800 6 wbs_dat_i[29]
port 337 nsew signal input
rlabel metal2 s 21362 0 21418 800 6 wbs_dat_i[2]
port 338 nsew signal input
rlabel metal2 s 140594 0 140650 800 6 wbs_dat_i[30]
port 339 nsew signal input
rlabel metal2 s 144734 0 144790 800 6 wbs_dat_i[31]
port 340 nsew signal input
rlabel metal2 s 26974 0 27030 800 6 wbs_dat_i[3]
port 341 nsew signal input
rlabel metal2 s 32494 0 32550 800 6 wbs_dat_i[4]
port 342 nsew signal input
rlabel metal2 s 36634 0 36690 800 6 wbs_dat_i[5]
port 343 nsew signal input
rlabel metal2 s 40774 0 40830 800 6 wbs_dat_i[6]
port 344 nsew signal input
rlabel metal2 s 45006 0 45062 800 6 wbs_dat_i[7]
port 345 nsew signal input
rlabel metal2 s 49146 0 49202 800 6 wbs_dat_i[8]
port 346 nsew signal input
rlabel metal2 s 53286 0 53342 800 6 wbs_dat_i[9]
port 347 nsew signal input
rlabel metal2 s 11702 0 11758 800 6 wbs_dat_o[0]
port 348 nsew signal output
rlabel metal2 s 58806 0 58862 800 6 wbs_dat_o[10]
port 349 nsew signal output
rlabel metal2 s 62946 0 63002 800 6 wbs_dat_o[11]
port 350 nsew signal output
rlabel metal2 s 67178 0 67234 800 6 wbs_dat_o[12]
port 351 nsew signal output
rlabel metal2 s 71318 0 71374 800 6 wbs_dat_o[13]
port 352 nsew signal output
rlabel metal2 s 75458 0 75514 800 6 wbs_dat_o[14]
port 353 nsew signal output
rlabel metal2 s 79598 0 79654 800 6 wbs_dat_o[15]
port 354 nsew signal output
rlabel metal2 s 83738 0 83794 800 6 wbs_dat_o[16]
port 355 nsew signal output
rlabel metal2 s 87878 0 87934 800 6 wbs_dat_o[17]
port 356 nsew signal output
rlabel metal2 s 92110 0 92166 800 6 wbs_dat_o[18]
port 357 nsew signal output
rlabel metal2 s 96250 0 96306 800 6 wbs_dat_o[19]
port 358 nsew signal output
rlabel metal2 s 17222 0 17278 800 6 wbs_dat_o[1]
port 359 nsew signal output
rlabel metal2 s 100390 0 100446 800 6 wbs_dat_o[20]
port 360 nsew signal output
rlabel metal2 s 104530 0 104586 800 6 wbs_dat_o[21]
port 361 nsew signal output
rlabel metal2 s 108670 0 108726 800 6 wbs_dat_o[22]
port 362 nsew signal output
rlabel metal2 s 112902 0 112958 800 6 wbs_dat_o[23]
port 363 nsew signal output
rlabel metal2 s 117042 0 117098 800 6 wbs_dat_o[24]
port 364 nsew signal output
rlabel metal2 s 121182 0 121238 800 6 wbs_dat_o[25]
port 365 nsew signal output
rlabel metal2 s 125322 0 125378 800 6 wbs_dat_o[26]
port 366 nsew signal output
rlabel metal2 s 129462 0 129518 800 6 wbs_dat_o[27]
port 367 nsew signal output
rlabel metal2 s 133694 0 133750 800 6 wbs_dat_o[28]
port 368 nsew signal output
rlabel metal2 s 137834 0 137890 800 6 wbs_dat_o[29]
port 369 nsew signal output
rlabel metal2 s 22834 0 22890 800 6 wbs_dat_o[2]
port 370 nsew signal output
rlabel metal2 s 141974 0 142030 800 6 wbs_dat_o[30]
port 371 nsew signal output
rlabel metal2 s 146114 0 146170 800 6 wbs_dat_o[31]
port 372 nsew signal output
rlabel metal2 s 28354 0 28410 800 6 wbs_dat_o[3]
port 373 nsew signal output
rlabel metal2 s 33874 0 33930 800 6 wbs_dat_o[4]
port 374 nsew signal output
rlabel metal2 s 38014 0 38070 800 6 wbs_dat_o[5]
port 375 nsew signal output
rlabel metal2 s 42154 0 42210 800 6 wbs_dat_o[6]
port 376 nsew signal output
rlabel metal2 s 46386 0 46442 800 6 wbs_dat_o[7]
port 377 nsew signal output
rlabel metal2 s 50526 0 50582 800 6 wbs_dat_o[8]
port 378 nsew signal output
rlabel metal2 s 54666 0 54722 800 6 wbs_dat_o[9]
port 379 nsew signal output
rlabel metal2 s 13082 0 13138 800 6 wbs_sel_i[0]
port 380 nsew signal input
rlabel metal2 s 18602 0 18658 800 6 wbs_sel_i[1]
port 381 nsew signal input
rlabel metal2 s 24214 0 24270 800 6 wbs_sel_i[2]
port 382 nsew signal input
rlabel metal2 s 29734 0 29790 800 6 wbs_sel_i[3]
port 383 nsew signal input
rlabel metal2 s 6182 0 6238 800 6 wbs_stb_i
port 384 nsew signal input
rlabel metal2 s 7562 0 7618 800 6 wbs_we_i
port 385 nsew signal input
<< properties >>
string LEFclass BLOCK
string FIXED_BBOX 0 0 198160 200304
string LEFview TRUE
string GDS_FILE /project/openlane/user_proj/runs/user_proj/results/magic/user_proj.gds
string GDS_END 98180260
string GDS_START 1540148
<< end >>

