magic
tech sky130A
magscale 1 2
timestamp 1645332165
<< locali >>
rect 215585 241927 215619 242641
rect 48881 239819 48915 239921
rect 43545 239479 43579 239717
rect 43637 239139 43671 239445
rect 49617 238935 49651 239717
rect 52377 238799 52411 239717
rect 54861 238867 54895 239717
rect 56241 239071 56275 239717
rect 57529 239003 57563 239717
rect 57713 238255 57747 239717
rect 59185 238323 59219 239717
rect 60105 239139 60139 239717
rect 62129 239479 62163 239717
rect 73445 238323 73479 239717
rect 75837 238255 75871 239717
rect 82921 239411 82955 239717
rect 97457 239411 97491 239717
rect 128829 239479 128863 239717
rect 168481 239275 168515 239649
rect 169309 239343 169343 239649
rect 171885 239547 171919 239921
rect 237941 239819 237975 239989
rect 177037 239207 177071 239649
rect 106933 3655 106967 3825
rect 117053 3723 117087 3825
<< viali >>
rect 215585 242641 215619 242675
rect 215585 241893 215619 241927
rect 237941 239989 237975 240023
rect 48881 239921 48915 239955
rect 48881 239785 48915 239819
rect 171885 239921 171919 239955
rect 43545 239717 43579 239751
rect 49617 239717 49651 239751
rect 43545 239445 43579 239479
rect 43637 239445 43671 239479
rect 43637 239105 43671 239139
rect 49617 238901 49651 238935
rect 52377 239717 52411 239751
rect 54861 239717 54895 239751
rect 56241 239717 56275 239751
rect 56241 239037 56275 239071
rect 57529 239717 57563 239751
rect 57529 238969 57563 239003
rect 57713 239717 57747 239751
rect 54861 238833 54895 238867
rect 52377 238765 52411 238799
rect 59185 239717 59219 239751
rect 60105 239717 60139 239751
rect 62129 239717 62163 239751
rect 62129 239445 62163 239479
rect 73445 239717 73479 239751
rect 60105 239105 60139 239139
rect 59185 238289 59219 238323
rect 73445 238289 73479 238323
rect 75837 239717 75871 239751
rect 57713 238221 57747 238255
rect 82921 239717 82955 239751
rect 82921 239377 82955 239411
rect 97457 239717 97491 239751
rect 128829 239717 128863 239751
rect 128829 239445 128863 239479
rect 168481 239649 168515 239683
rect 97457 239377 97491 239411
rect 169309 239649 169343 239683
rect 237941 239785 237975 239819
rect 171885 239513 171919 239547
rect 177037 239649 177071 239683
rect 169309 239309 169343 239343
rect 168481 239241 168515 239275
rect 177037 239173 177071 239207
rect 75837 238221 75871 238255
rect 106933 3825 106967 3859
rect 117053 3825 117087 3859
rect 117053 3689 117087 3723
rect 106933 3621 106967 3655
<< metal1 >>
rect 201494 702992 201500 703044
rect 201552 703032 201558 703044
rect 202782 703032 202788 703044
rect 201552 703004 202788 703032
rect 201552 702992 201558 703004
rect 202782 702992 202788 703004
rect 202840 702992 202846 703044
rect 229738 700952 229744 701004
rect 229796 700992 229802 701004
rect 267642 700992 267648 701004
rect 229796 700964 267648 700992
rect 229796 700952 229802 700964
rect 267642 700952 267648 700964
rect 267700 700952 267706 701004
rect 211798 700884 211804 700936
rect 211856 700924 211862 700936
rect 332502 700924 332508 700936
rect 211856 700896 332508 700924
rect 211856 700884 211862 700896
rect 332502 700884 332508 700896
rect 332560 700884 332566 700936
rect 220078 700816 220084 700868
rect 220136 700856 220142 700868
rect 348786 700856 348792 700868
rect 220136 700828 348792 700856
rect 220136 700816 220142 700828
rect 348786 700816 348792 700828
rect 348844 700816 348850 700868
rect 193858 700748 193864 700800
rect 193916 700788 193922 700800
rect 364978 700788 364984 700800
rect 193916 700760 364984 700788
rect 193916 700748 193922 700760
rect 364978 700748 364984 700760
rect 365036 700748 365042 700800
rect 209038 700680 209044 700732
rect 209096 700720 209102 700732
rect 397454 700720 397460 700732
rect 209096 700692 397460 700720
rect 209096 700680 209102 700692
rect 397454 700680 397460 700692
rect 397512 700680 397518 700732
rect 215938 700612 215944 700664
rect 215996 700652 216002 700664
rect 413646 700652 413652 700664
rect 215996 700624 413652 700652
rect 215996 700612 216002 700624
rect 413646 700612 413652 700624
rect 413704 700612 413710 700664
rect 191098 700544 191104 700596
rect 191156 700584 191162 700596
rect 429838 700584 429844 700596
rect 191156 700556 429844 700584
rect 191156 700544 191162 700556
rect 429838 700544 429844 700556
rect 429896 700544 429902 700596
rect 204898 700476 204904 700528
rect 204956 700516 204962 700528
rect 462314 700516 462320 700528
rect 204956 700488 462320 700516
rect 204956 700476 204962 700488
rect 462314 700476 462320 700488
rect 462372 700476 462378 700528
rect 170306 700408 170312 700460
rect 170364 700448 170370 700460
rect 176838 700448 176844 700460
rect 170364 700420 176844 700448
rect 170364 700408 170370 700420
rect 176838 700408 176844 700420
rect 176896 700408 176902 700460
rect 197998 700408 198004 700460
rect 198056 700448 198062 700460
rect 235166 700448 235172 700460
rect 198056 700420 235172 700448
rect 198056 700408 198062 700420
rect 235166 700408 235172 700420
rect 235224 700408 235230 700460
rect 238018 700408 238024 700460
rect 238076 700448 238082 700460
rect 527174 700448 527180 700460
rect 238076 700420 527180 700448
rect 238076 700408 238082 700420
rect 527174 700408 527180 700420
rect 527232 700408 527238 700460
rect 137830 700340 137836 700392
rect 137888 700380 137894 700392
rect 176746 700380 176752 700392
rect 137888 700352 176752 700380
rect 137888 700340 137894 700352
rect 176746 700340 176752 700352
rect 176804 700340 176810 700392
rect 189718 700340 189724 700392
rect 189776 700380 189782 700392
rect 494790 700380 494796 700392
rect 189776 700352 494796 700380
rect 189776 700340 189782 700352
rect 494790 700340 494796 700352
rect 494848 700340 494854 700392
rect 89162 700272 89168 700324
rect 89220 700312 89226 700324
rect 176654 700312 176660 700324
rect 89220 700284 176660 700312
rect 89220 700272 89226 700284
rect 176654 700272 176660 700284
rect 176712 700272 176718 700324
rect 185578 700272 185584 700324
rect 185636 700312 185642 700324
rect 559650 700312 559656 700324
rect 185636 700284 559656 700312
rect 185636 700272 185642 700284
rect 559650 700272 559656 700284
rect 559708 700272 559714 700324
rect 24302 699660 24308 699712
rect 24360 699700 24366 699712
rect 24762 699700 24768 699712
rect 24360 699672 24768 699700
rect 24360 699660 24366 699672
rect 24762 699660 24768 699672
rect 24820 699660 24826 699712
rect 39850 699660 39856 699712
rect 39908 699700 39914 699712
rect 40494 699700 40500 699712
rect 39908 699672 40500 699700
rect 39908 699660 39914 699672
rect 40494 699660 40500 699672
rect 40552 699660 40558 699712
rect 71774 699660 71780 699712
rect 71832 699700 71838 699712
rect 72970 699700 72976 699712
rect 71832 699672 72976 699700
rect 71832 699660 71838 699672
rect 72970 699660 72976 699672
rect 73028 699660 73034 699712
rect 105446 699660 105452 699712
rect 105504 699700 105510 699712
rect 106182 699700 106188 699712
rect 105504 699672 106188 699700
rect 105504 699660 105510 699672
rect 106182 699660 106188 699672
rect 106240 699660 106246 699712
rect 196618 696940 196624 696992
rect 196676 696980 196682 696992
rect 580166 696980 580172 696992
rect 196676 696952 580172 696980
rect 196676 696940 196682 696952
rect 580166 696940 580172 696952
rect 580224 696940 580230 696992
rect 2774 683612 2780 683664
rect 2832 683652 2838 683664
rect 6178 683652 6184 683664
rect 2832 683624 6184 683652
rect 2832 683612 2838 683624
rect 6178 683612 6184 683624
rect 6236 683612 6242 683664
rect 182818 670692 182824 670744
rect 182876 670732 182882 670744
rect 580166 670732 580172 670744
rect 182876 670704 580172 670732
rect 182876 670692 182882 670704
rect 580166 670692 580172 670704
rect 580224 670692 580230 670744
rect 3510 656888 3516 656940
rect 3568 656928 3574 656940
rect 21358 656928 21364 656940
rect 3568 656900 21364 656928
rect 3568 656888 3574 656900
rect 21358 656888 21364 656900
rect 21416 656888 21422 656940
rect 200758 643084 200764 643136
rect 200816 643124 200822 643136
rect 580166 643124 580172 643136
rect 200816 643096 580172 643124
rect 200816 643084 200822 643096
rect 580166 643084 580172 643096
rect 580224 643084 580230 643136
rect 3510 632068 3516 632120
rect 3568 632108 3574 632120
rect 15838 632108 15844 632120
rect 3568 632080 15844 632108
rect 3568 632068 3574 632080
rect 15838 632068 15844 632080
rect 15896 632068 15902 632120
rect 214558 630640 214564 630692
rect 214616 630680 214622 630692
rect 579982 630680 579988 630692
rect 214616 630652 579988 630680
rect 214616 630640 214622 630652
rect 579982 630640 579988 630652
rect 580040 630640 580046 630692
rect 180058 616836 180064 616888
rect 180116 616876 180122 616888
rect 580166 616876 580172 616888
rect 180116 616848 580172 616876
rect 180116 616836 180122 616848
rect 580166 616836 580172 616848
rect 580224 616836 580230 616888
rect 3326 605820 3332 605872
rect 3384 605860 3390 605872
rect 25498 605860 25504 605872
rect 3384 605832 25504 605860
rect 3384 605820 3390 605832
rect 25498 605820 25504 605832
rect 25556 605820 25562 605872
rect 226978 590656 226984 590708
rect 227036 590696 227042 590708
rect 580166 590696 580172 590708
rect 227036 590668 580172 590696
rect 227036 590656 227042 590668
rect 580166 590656 580172 590668
rect 580224 590656 580230 590708
rect 3326 579640 3332 579692
rect 3384 579680 3390 579692
rect 10318 579680 10324 579692
rect 3384 579652 10324 579680
rect 3384 579640 3390 579652
rect 10318 579640 10324 579652
rect 10376 579640 10382 579692
rect 231118 563048 231124 563100
rect 231176 563088 231182 563100
rect 579890 563088 579896 563100
rect 231176 563060 579896 563088
rect 231176 563048 231182 563060
rect 579890 563048 579896 563060
rect 579948 563048 579954 563100
rect 3326 553392 3332 553444
rect 3384 553432 3390 553444
rect 28258 553432 28264 553444
rect 3384 553404 28264 553432
rect 3384 553392 3390 553404
rect 28258 553392 28264 553404
rect 28316 553392 28322 553444
rect 269758 536800 269764 536852
rect 269816 536840 269822 536852
rect 580166 536840 580172 536852
rect 269816 536812 580172 536840
rect 269816 536800 269822 536812
rect 580166 536800 580172 536812
rect 580224 536800 580230 536852
rect 3326 527144 3332 527196
rect 3384 527184 3390 527196
rect 13078 527184 13084 527196
rect 3384 527156 13084 527184
rect 3384 527144 3390 527156
rect 13078 527144 13084 527156
rect 13136 527144 13142 527196
rect 266998 524424 267004 524476
rect 267056 524464 267062 524476
rect 580166 524464 580172 524476
rect 267056 524436 580172 524464
rect 267056 524424 267062 524436
rect 580166 524424 580172 524436
rect 580224 524424 580230 524476
rect 3326 514768 3332 514820
rect 3384 514808 3390 514820
rect 35158 514808 35164 514820
rect 3384 514780 35164 514808
rect 3384 514768 3390 514780
rect 35158 514768 35164 514780
rect 35216 514768 35222 514820
rect 265618 510620 265624 510672
rect 265676 510660 265682 510672
rect 580166 510660 580172 510672
rect 265676 510632 580172 510660
rect 265676 510620 265682 510632
rect 580166 510620 580172 510632
rect 580224 510620 580230 510672
rect 2866 500964 2872 501016
rect 2924 501004 2930 501016
rect 31018 501004 31024 501016
rect 2924 500976 31024 501004
rect 2924 500964 2930 500976
rect 31018 500964 31024 500976
rect 31076 500964 31082 501016
rect 268378 484372 268384 484424
rect 268436 484412 268442 484424
rect 580166 484412 580172 484424
rect 268436 484384 580172 484412
rect 268436 484372 268442 484384
rect 580166 484372 580172 484384
rect 580224 484372 580230 484424
rect 3326 474716 3332 474768
rect 3384 474756 3390 474768
rect 14458 474756 14464 474768
rect 3384 474728 14464 474756
rect 3384 474716 3390 474728
rect 14458 474716 14464 474728
rect 14516 474716 14522 474768
rect 153194 472608 153200 472660
rect 153252 472648 153258 472660
rect 176930 472648 176936 472660
rect 153252 472620 176936 472648
rect 153252 472608 153258 472620
rect 176930 472608 176936 472620
rect 176988 472608 176994 472660
rect 3326 462340 3332 462392
rect 3384 462380 3390 462392
rect 19978 462380 19984 462392
rect 3384 462352 19984 462380
rect 3384 462340 3390 462352
rect 19978 462340 19984 462352
rect 20036 462340 20042 462392
rect 479518 456764 479524 456816
rect 479576 456804 479582 456816
rect 579614 456804 579620 456816
rect 479576 456776 579620 456804
rect 479576 456764 479582 456776
rect 579614 456764 579620 456776
rect 579672 456764 579678 456816
rect 3326 448536 3332 448588
rect 3384 448576 3390 448588
rect 32398 448576 32404 448588
rect 3384 448548 32404 448576
rect 3384 448536 3390 448548
rect 32398 448536 32404 448548
rect 32456 448536 32462 448588
rect 39758 425688 39764 425740
rect 39816 425728 39822 425740
rect 71774 425728 71780 425740
rect 39816 425700 71780 425728
rect 39816 425688 39822 425700
rect 71774 425688 71780 425700
rect 71832 425688 71838 425740
rect 106182 425688 106188 425740
rect 106240 425728 106246 425740
rect 177022 425728 177028 425740
rect 106240 425700 177028 425728
rect 106240 425688 106246 425700
rect 177022 425688 177028 425700
rect 177080 425688 177086 425740
rect 3142 422288 3148 422340
rect 3200 422328 3206 422340
rect 17218 422328 17224 422340
rect 3200 422300 17224 422328
rect 3200 422288 3206 422300
rect 17218 422288 17224 422300
rect 17276 422288 17282 422340
rect 486418 418140 486424 418192
rect 486476 418180 486482 418192
rect 579706 418180 579712 418192
rect 486476 418152 579712 418180
rect 486476 418140 486482 418152
rect 579706 418140 579712 418152
rect 579764 418140 579770 418192
rect 482278 404336 482284 404388
rect 482336 404376 482342 404388
rect 580166 404376 580172 404388
rect 482336 404348 580172 404376
rect 482336 404336 482342 404348
rect 580166 404336 580172 404348
rect 580224 404336 580230 404388
rect 3326 397468 3332 397520
rect 3384 397508 3390 397520
rect 33778 397508 33784 397520
rect 3384 397480 33784 397508
rect 3384 397468 3390 397480
rect 33778 397468 33784 397480
rect 33836 397468 33842 397520
rect 483658 378156 483664 378208
rect 483716 378196 483722 378208
rect 580166 378196 580172 378208
rect 483716 378168 580172 378196
rect 483716 378156 483722 378168
rect 580166 378156 580172 378168
rect 580224 378156 580230 378208
rect 294598 376728 294604 376780
rect 294656 376768 294662 376780
rect 337654 376768 337660 376780
rect 294656 376740 337660 376768
rect 294656 376728 294662 376740
rect 337654 376728 337660 376740
rect 337712 376728 337718 376780
rect 262858 375368 262864 375420
rect 262916 375408 262922 375420
rect 337746 375408 337752 375420
rect 262916 375380 337752 375408
rect 262916 375368 262922 375380
rect 337746 375368 337752 375380
rect 337804 375368 337810 375420
rect 291838 372580 291844 372632
rect 291896 372620 291902 372632
rect 337470 372620 337476 372632
rect 291896 372592 337476 372620
rect 291896 372580 291902 372592
rect 337470 372580 337476 372592
rect 337528 372580 337534 372632
rect 3326 371220 3332 371272
rect 3384 371260 3390 371272
rect 20070 371260 20076 371272
rect 3384 371232 20076 371260
rect 3384 371220 3390 371232
rect 20070 371220 20076 371232
rect 20128 371220 20134 371272
rect 261478 369928 261484 369980
rect 261536 369968 261542 369980
rect 337470 369968 337476 369980
rect 261536 369940 337476 369968
rect 261536 369928 261542 369940
rect 337470 369928 337476 369940
rect 337528 369928 337534 369980
rect 35618 369860 35624 369912
rect 35676 369900 35682 369912
rect 37918 369900 37924 369912
rect 35676 369872 37924 369900
rect 35676 369860 35682 369872
rect 37918 369860 37924 369872
rect 37976 369860 37982 369912
rect 258718 369860 258724 369912
rect 258776 369900 258782 369912
rect 337746 369900 337752 369912
rect 258776 369872 337752 369900
rect 258776 369860 258782 369872
rect 337746 369860 337752 369872
rect 337804 369860 337810 369912
rect 195882 367072 195888 367124
rect 195940 367112 195946 367124
rect 337470 367112 337476 367124
rect 195940 367084 337476 367112
rect 195940 367072 195946 367084
rect 337470 367072 337476 367084
rect 337528 367072 337534 367124
rect 485038 364352 485044 364404
rect 485096 364392 485102 364404
rect 580166 364392 580172 364404
rect 485096 364364 580172 364392
rect 485096 364352 485102 364364
rect 580166 364352 580172 364364
rect 580224 364352 580230 364404
rect 480898 351908 480904 351960
rect 480956 351948 480962 351960
rect 580166 351948 580172 351960
rect 480956 351920 580172 351948
rect 480956 351908 480962 351920
rect 580166 351908 580172 351920
rect 580224 351908 580230 351960
rect 187602 349120 187608 349172
rect 187660 349160 187666 349172
rect 337746 349160 337752 349172
rect 187660 349132 337752 349160
rect 187660 349120 187666 349132
rect 337746 349120 337752 349132
rect 337804 349120 337810 349172
rect 35802 347828 35808 347880
rect 35860 347868 35866 347880
rect 37642 347868 37648 347880
rect 35860 347840 37648 347868
rect 35860 347828 35866 347840
rect 37642 347828 37648 347840
rect 37700 347828 37706 347880
rect 254578 347760 254584 347812
rect 254636 347800 254642 347812
rect 337654 347800 337660 347812
rect 254636 347772 337660 347800
rect 254636 347760 254642 347772
rect 337654 347760 337660 347772
rect 337712 347760 337718 347812
rect 3050 345040 3056 345092
rect 3108 345080 3114 345092
rect 35250 345080 35256 345092
rect 3108 345052 35256 345080
rect 3108 345040 3114 345052
rect 35250 345040 35256 345052
rect 35308 345040 35314 345092
rect 35158 339396 35164 339448
rect 35216 339436 35222 339448
rect 146294 339436 146300 339448
rect 35216 339408 146300 339436
rect 35216 339396 35222 339408
rect 146294 339396 146300 339408
rect 146352 339396 146358 339448
rect 3418 339328 3424 339380
rect 3476 339368 3482 339380
rect 133874 339368 133880 339380
rect 3476 339340 133880 339368
rect 3476 339328 3482 339340
rect 133874 339328 133880 339340
rect 133932 339328 133938 339380
rect 3510 339260 3516 339312
rect 3568 339300 3574 339312
rect 138014 339300 138020 339312
rect 3568 339272 138020 339300
rect 3568 339260 3574 339272
rect 138014 339260 138020 339272
rect 138072 339260 138078 339312
rect 100662 339192 100668 339244
rect 100720 339232 100726 339244
rect 238018 339232 238024 339244
rect 100720 339204 238024 339232
rect 100720 339192 100726 339204
rect 238018 339192 238024 339204
rect 238076 339192 238082 339244
rect 3602 339124 3608 339176
rect 3660 339164 3666 339176
rect 142154 339164 142160 339176
rect 3660 339136 142160 339164
rect 3660 339124 3666 339136
rect 142154 339124 142160 339136
rect 142212 339124 142218 339176
rect 3786 339056 3792 339108
rect 3844 339096 3850 339108
rect 157334 339096 157340 339108
rect 3844 339068 157340 339096
rect 3844 339056 3850 339068
rect 157334 339056 157340 339068
rect 157392 339056 157398 339108
rect 38746 338988 38752 339040
rect 38804 339028 38810 339040
rect 202966 339028 202972 339040
rect 38804 339000 202972 339028
rect 38804 338988 38810 339000
rect 202966 338988 202972 339000
rect 203024 338988 203030 339040
rect 38378 338920 38384 338972
rect 38436 338960 38442 338972
rect 240686 338960 240692 338972
rect 38436 338932 240692 338960
rect 38436 338920 38442 338932
rect 240686 338920 240692 338932
rect 240744 338920 240750 338972
rect 97902 338852 97908 338904
rect 97960 338892 97966 338904
rect 580258 338892 580264 338904
rect 97960 338864 580264 338892
rect 97960 338852 97966 338864
rect 580258 338852 580264 338864
rect 580316 338852 580322 338904
rect 89530 338784 89536 338836
rect 89588 338824 89594 338836
rect 580350 338824 580356 338836
rect 89588 338796 580356 338824
rect 89588 338784 89594 338796
rect 580350 338784 580356 338796
rect 580408 338784 580414 338836
rect 82722 338716 82728 338768
rect 82780 338756 82786 338768
rect 580534 338756 580540 338768
rect 82780 338728 580540 338756
rect 82780 338716 82786 338728
rect 580534 338716 580540 338728
rect 580592 338716 580598 338768
rect 39850 338648 39856 338700
rect 39908 338688 39914 338700
rect 128354 338688 128360 338700
rect 39908 338660 128360 338688
rect 39908 338648 39914 338660
rect 128354 338648 128360 338660
rect 128412 338648 128418 338700
rect 121362 338580 121368 338632
rect 121420 338620 121426 338632
rect 176838 338620 176844 338632
rect 121420 338592 176844 338620
rect 121420 338580 121426 338592
rect 176838 338580 176844 338592
rect 176896 338580 176902 338632
rect 38562 338036 38568 338088
rect 38620 338076 38626 338088
rect 337378 338076 337384 338088
rect 38620 338048 337384 338076
rect 38620 338036 38626 338048
rect 337378 338036 337384 338048
rect 337436 338036 337442 338088
rect 42058 337832 42064 337884
rect 42116 337872 42122 337884
rect 379514 337872 379520 337884
rect 42116 337844 379520 337872
rect 42116 337832 42122 337844
rect 379514 337832 379520 337844
rect 379572 337832 379578 337884
rect 50338 337764 50344 337816
rect 50396 337804 50402 337816
rect 394694 337804 394700 337816
rect 50396 337776 394700 337804
rect 50396 337764 50402 337776
rect 394694 337764 394700 337776
rect 394752 337764 394758 337816
rect 78582 337696 78588 337748
rect 78640 337736 78646 337748
rect 78640 337708 84194 337736
rect 78640 337696 78646 337708
rect 56502 337628 56508 337680
rect 56560 337668 56566 337680
rect 61378 337668 61384 337680
rect 56560 337640 61384 337668
rect 56560 337628 56566 337640
rect 61378 337628 61384 337640
rect 61436 337628 61442 337680
rect 77202 337628 77208 337680
rect 77260 337668 77266 337680
rect 79318 337668 79324 337680
rect 77260 337640 79324 337668
rect 77260 337628 77266 337640
rect 79318 337628 79324 337640
rect 79376 337628 79382 337680
rect 84166 337668 84194 337708
rect 122742 337696 122748 337748
rect 122800 337736 122806 337748
rect 176746 337736 176752 337748
rect 122800 337708 176752 337736
rect 122800 337696 122806 337708
rect 176746 337696 176752 337708
rect 176804 337696 176810 337748
rect 388438 337696 388444 337748
rect 388496 337736 388502 337748
rect 391934 337736 391940 337748
rect 388496 337708 391940 337736
rect 388496 337696 388502 337708
rect 391934 337696 391940 337708
rect 391992 337696 391998 337748
rect 126238 337668 126244 337680
rect 84166 337640 126244 337668
rect 126238 337628 126244 337640
rect 126296 337628 126302 337680
rect 143442 337628 143448 337680
rect 143500 337668 143506 337680
rect 241514 337668 241520 337680
rect 143500 337640 241520 337668
rect 143500 337628 143506 337640
rect 241514 337628 241520 337640
rect 241572 337628 241578 337680
rect 367738 337628 367744 337680
rect 367796 337668 367802 337680
rect 369854 337668 369860 337680
rect 367796 337640 369860 337668
rect 367796 337628 367802 337640
rect 369854 337628 369860 337640
rect 369912 337628 369918 337680
rect 387058 337628 387064 337680
rect 387116 337668 387122 337680
rect 389174 337668 389180 337680
rect 387116 337640 389180 337668
rect 387116 337628 387122 337640
rect 389174 337628 389180 337640
rect 389232 337628 389238 337680
rect 118602 337560 118608 337612
rect 118660 337600 118666 337612
rect 237742 337600 237748 337612
rect 118660 337572 237748 337600
rect 118660 337560 118666 337572
rect 237742 337560 237748 337572
rect 237800 337560 237806 337612
rect 117222 337492 117228 337544
rect 117280 337532 117286 337544
rect 237650 337532 237656 337544
rect 117280 337504 237656 337532
rect 117280 337492 117286 337504
rect 237650 337492 237656 337504
rect 237708 337492 237714 337544
rect 355318 337492 355324 337544
rect 355376 337532 355382 337544
rect 372614 337532 372620 337544
rect 355376 337504 372620 337532
rect 355376 337492 355382 337504
rect 372614 337492 372620 337504
rect 372672 337492 372678 337544
rect 104802 337424 104808 337476
rect 104860 337464 104866 337476
rect 237558 337464 237564 337476
rect 104860 337436 237564 337464
rect 104860 337424 104866 337436
rect 237558 337424 237564 337436
rect 237616 337424 237622 337476
rect 364978 337424 364984 337476
rect 365036 337464 365042 337476
rect 397454 337464 397460 337476
rect 365036 337436 397460 337464
rect 365036 337424 365042 337436
rect 397454 337424 397460 337436
rect 397512 337424 397518 337476
rect 43438 337356 43444 337408
rect 43496 337396 43502 337408
rect 96614 337396 96620 337408
rect 43496 337368 96620 337396
rect 43496 337356 43502 337368
rect 96614 337356 96620 337368
rect 96672 337356 96678 337408
rect 99282 337356 99288 337408
rect 99340 337396 99346 337408
rect 236638 337396 236644 337408
rect 99340 337368 236644 337396
rect 99340 337356 99346 337368
rect 236638 337356 236644 337368
rect 236696 337356 236702 337408
rect 349798 337356 349804 337408
rect 349856 337396 349862 337408
rect 385034 337396 385040 337408
rect 349856 337368 385040 337396
rect 349856 337356 349862 337368
rect 385034 337356 385040 337368
rect 385092 337356 385098 337408
rect 387794 337396 387800 337408
rect 385512 337368 387800 337396
rect 93578 337288 93584 337340
rect 93636 337328 93642 337340
rect 232498 337328 232504 337340
rect 93636 337300 232504 337328
rect 93636 337288 93642 337300
rect 232498 337288 232504 337300
rect 232556 337288 232562 337340
rect 352558 337288 352564 337340
rect 352616 337328 352622 337340
rect 385512 337328 385540 337368
rect 387794 337356 387800 337368
rect 387852 337356 387858 337408
rect 352616 337300 385540 337328
rect 352616 337288 352622 337300
rect 385678 337288 385684 337340
rect 385736 337328 385742 337340
rect 390554 337328 390560 337340
rect 385736 337300 390560 337328
rect 385736 337288 385742 337300
rect 390554 337288 390560 337300
rect 390612 337288 390618 337340
rect 89622 337220 89628 337272
rect 89680 337260 89686 337272
rect 238294 337260 238300 337272
rect 89680 337232 238300 337260
rect 89680 337220 89686 337232
rect 238294 337220 238300 337232
rect 238352 337220 238358 337272
rect 287698 337220 287704 337272
rect 287756 337260 287762 337272
rect 382274 337260 382280 337272
rect 287756 337232 382280 337260
rect 287756 337220 287762 337232
rect 382274 337220 382280 337232
rect 382332 337220 382338 337272
rect 84010 337152 84016 337204
rect 84068 337192 84074 337204
rect 238202 337192 238208 337204
rect 84068 337164 238208 337192
rect 84068 337152 84074 337164
rect 238202 337152 238208 337164
rect 238260 337152 238266 337204
rect 255958 337152 255964 337204
rect 256016 337192 256022 337204
rect 371234 337192 371240 337204
rect 256016 337164 371240 337192
rect 256016 337152 256022 337164
rect 371234 337152 371240 337164
rect 371292 337152 371298 337204
rect 382918 337152 382924 337204
rect 382976 337192 382982 337204
rect 386414 337192 386420 337204
rect 382976 337164 386420 337192
rect 382976 337152 382982 337164
rect 386414 337152 386420 337164
rect 386472 337152 386478 337204
rect 40494 337084 40500 337136
rect 40552 337124 40558 337136
rect 60734 337124 60740 337136
rect 40552 337096 60740 337124
rect 40552 337084 40558 337096
rect 60734 337084 60740 337096
rect 60792 337084 60798 337136
rect 67542 337084 67548 337136
rect 67600 337124 67606 337136
rect 236730 337124 236736 337136
rect 67600 337096 236736 337124
rect 67600 337084 67606 337096
rect 236730 337084 236736 337096
rect 236788 337084 236794 337136
rect 249058 337084 249064 337136
rect 249116 337124 249122 337136
rect 375374 337124 375380 337136
rect 249116 337096 375380 337124
rect 249116 337084 249122 337096
rect 375374 337084 375380 337096
rect 375432 337084 375438 337136
rect 381538 337084 381544 337136
rect 381596 337124 381602 337136
rect 386506 337124 386512 337136
rect 381596 337096 386512 337124
rect 381596 337084 381602 337096
rect 386506 337084 386512 337096
rect 386564 337084 386570 337136
rect 38378 337016 38384 337068
rect 38436 337056 38442 337068
rect 59354 337056 59360 337068
rect 38436 337028 59360 337056
rect 38436 337016 38442 337028
rect 59354 337016 59360 337028
rect 59412 337016 59418 337068
rect 66162 337016 66168 337068
rect 66220 337056 66226 337068
rect 239398 337056 239404 337068
rect 66220 337028 239404 337056
rect 66220 337016 66226 337028
rect 239398 337016 239404 337028
rect 239456 337016 239462 337068
rect 251818 337016 251824 337068
rect 251876 337056 251882 337068
rect 433334 337056 433340 337068
rect 251876 337028 433340 337056
rect 251876 337016 251882 337028
rect 433334 337016 433340 337028
rect 433392 337016 433398 337068
rect 46198 336948 46204 337000
rect 46256 336988 46262 337000
rect 379422 336988 379428 337000
rect 46256 336960 379428 336988
rect 46256 336948 46262 336960
rect 379422 336948 379428 336960
rect 379480 336948 379486 337000
rect 379514 336948 379520 337000
rect 379572 336988 379578 337000
rect 387794 336988 387800 337000
rect 379572 336960 387800 336988
rect 379572 336948 379578 336960
rect 387794 336948 387800 336960
rect 387852 336948 387858 337000
rect 411898 336948 411904 337000
rect 411956 336988 411962 337000
rect 440234 336988 440240 337000
rect 411956 336960 440240 336988
rect 411956 336948 411962 336960
rect 440234 336948 440240 336960
rect 440292 336948 440298 337000
rect 48958 336880 48964 336932
rect 49016 336920 49022 336932
rect 383746 336920 383752 336932
rect 49016 336892 383752 336920
rect 49016 336880 49022 336892
rect 383746 336880 383752 336892
rect 383804 336880 383810 336932
rect 402238 336880 402244 336932
rect 402296 336920 402302 336932
rect 407114 336920 407120 336932
rect 402296 336892 407120 336920
rect 402296 336880 402302 336892
rect 407114 336880 407120 336892
rect 407172 336880 407178 336932
rect 409138 336880 409144 336932
rect 409196 336920 409202 336932
rect 425054 336920 425060 336932
rect 409196 336892 425060 336920
rect 409196 336880 409202 336892
rect 425054 336880 425060 336892
rect 425112 336880 425118 336932
rect 384942 336812 384948 336864
rect 385000 336852 385006 336864
rect 396074 336852 396080 336864
rect 385000 336824 396080 336852
rect 385000 336812 385006 336824
rect 396074 336812 396080 336824
rect 396132 336812 396138 336864
rect 399478 336812 399484 336864
rect 399536 336852 399542 336864
rect 405734 336852 405740 336864
rect 399536 336824 405740 336852
rect 399536 336812 399542 336824
rect 405734 336812 405740 336824
rect 405792 336812 405798 336864
rect 406378 336812 406384 336864
rect 406436 336852 406442 336864
rect 422938 336852 422944 336864
rect 406436 336824 422944 336852
rect 406436 336812 406442 336824
rect 422938 336812 422944 336824
rect 422996 336812 423002 336864
rect 40310 336744 40316 336796
rect 40368 336784 40374 336796
rect 57974 336784 57980 336796
rect 40368 336756 57980 336784
rect 40368 336744 40374 336756
rect 57974 336744 57980 336756
rect 58032 336744 58038 336796
rect 70302 336744 70308 336796
rect 70360 336784 70366 336796
rect 75178 336784 75184 336796
rect 70360 336756 75184 336784
rect 70360 336744 70366 336756
rect 75178 336744 75184 336756
rect 75236 336744 75242 336796
rect 95142 336744 95148 336796
rect 95200 336784 95206 336796
rect 106918 336784 106924 336796
rect 95200 336756 106924 336784
rect 95200 336744 95206 336756
rect 106918 336744 106924 336756
rect 106976 336744 106982 336796
rect 351178 336744 351184 336796
rect 351236 336784 351242 336796
rect 364518 336784 364524 336796
rect 351236 336756 364524 336784
rect 351236 336744 351242 336756
rect 364518 336744 364524 336756
rect 364576 336744 364582 336796
rect 373258 336744 373264 336796
rect 373316 336784 373322 336796
rect 378134 336784 378140 336796
rect 373316 336756 378140 336784
rect 373316 336744 373322 336756
rect 378134 336744 378140 336756
rect 378192 336744 378198 336796
rect 391198 336744 391204 336796
rect 391256 336784 391262 336796
rect 393314 336784 393320 336796
rect 391256 336756 393320 336784
rect 391256 336744 391262 336756
rect 393314 336744 393320 336756
rect 393372 336744 393378 336796
rect 290458 336608 290464 336660
rect 290516 336648 290522 336660
rect 390554 336648 390560 336660
rect 290516 336620 390560 336648
rect 290516 336608 290522 336620
rect 390554 336608 390560 336620
rect 390612 336608 390618 336660
rect 81342 336540 81348 336592
rect 81400 336580 81406 336592
rect 173158 336580 173164 336592
rect 81400 336552 173164 336580
rect 81400 336540 81406 336552
rect 173158 336540 173164 336552
rect 173216 336540 173222 336592
rect 250438 336540 250444 336592
rect 250496 336580 250502 336592
rect 376846 336580 376852 336592
rect 250496 336552 376852 336580
rect 250496 336540 250502 336552
rect 376846 336540 376852 336552
rect 376904 336540 376910 336592
rect 131022 336472 131028 336524
rect 131080 336512 131086 336524
rect 225598 336512 225604 336524
rect 131080 336484 225604 336512
rect 131080 336472 131086 336484
rect 225598 336472 225604 336484
rect 225656 336472 225662 336524
rect 234522 336472 234528 336524
rect 234580 336512 234586 336524
rect 384942 336512 384948 336524
rect 234580 336484 384948 336512
rect 234580 336472 234586 336484
rect 384942 336472 384948 336484
rect 385000 336472 385006 336524
rect 129642 336404 129648 336456
rect 129700 336444 129706 336456
rect 175918 336444 175924 336456
rect 129700 336416 175924 336444
rect 129700 336404 129706 336416
rect 175918 336404 175924 336416
rect 175976 336404 175982 336456
rect 223482 336404 223488 336456
rect 223540 336444 223546 336456
rect 379514 336444 379520 336456
rect 223540 336416 379520 336444
rect 223540 336404 223546 336416
rect 379514 336404 379520 336416
rect 379572 336404 379578 336456
rect 81250 336336 81256 336388
rect 81308 336376 81314 336388
rect 177298 336376 177304 336388
rect 81308 336348 177304 336376
rect 81308 336336 81314 336348
rect 177298 336336 177304 336348
rect 177356 336336 177362 336388
rect 243538 336336 243544 336388
rect 243596 336376 243602 336388
rect 403250 336376 403256 336388
rect 243596 336348 403256 336376
rect 243596 336336 243602 336348
rect 403250 336336 403256 336348
rect 403308 336336 403314 336388
rect 37090 336268 37096 336320
rect 37148 336308 37154 336320
rect 97994 336308 98000 336320
rect 37148 336280 98000 336308
rect 37148 336268 37154 336280
rect 97994 336268 98000 336280
rect 98052 336268 98058 336320
rect 121270 336268 121276 336320
rect 121328 336308 121334 336320
rect 220814 336308 220820 336320
rect 121328 336280 220820 336308
rect 121328 336268 121334 336280
rect 220814 336268 220820 336280
rect 220872 336268 220878 336320
rect 244918 336268 244924 336320
rect 244976 336308 244982 336320
rect 409874 336308 409880 336320
rect 244976 336280 409880 336308
rect 244976 336268 244982 336280
rect 409874 336268 409880 336280
rect 409932 336268 409938 336320
rect 37182 336200 37188 336252
rect 37240 336240 37246 336252
rect 75914 336240 75920 336252
rect 37240 336212 75920 336240
rect 37240 336200 37246 336212
rect 75914 336200 75920 336212
rect 75972 336200 75978 336252
rect 96522 336200 96528 336252
rect 96580 336240 96586 336252
rect 207658 336240 207664 336252
rect 96580 336212 207664 336240
rect 96580 336200 96586 336212
rect 207658 336200 207664 336212
rect 207716 336200 207722 336252
rect 213822 336200 213828 336252
rect 213880 336240 213886 336252
rect 397454 336240 397460 336252
rect 213880 336212 397460 336240
rect 213880 336200 213886 336212
rect 397454 336200 397460 336212
rect 397512 336200 397518 336252
rect 19978 336132 19984 336184
rect 20036 336172 20042 336184
rect 150434 336172 150440 336184
rect 20036 336144 150440 336172
rect 20036 336132 20042 336144
rect 150434 336132 150440 336144
rect 150492 336132 150498 336184
rect 247678 336132 247684 336184
rect 247736 336172 247742 336184
rect 442994 336172 443000 336184
rect 247736 336144 443000 336172
rect 247736 336132 247742 336144
rect 442994 336132 443000 336144
rect 443052 336132 443058 336184
rect 35710 336064 35716 336116
rect 35768 336104 35774 336116
rect 371234 336104 371240 336116
rect 35768 336076 371240 336104
rect 35768 336064 35774 336076
rect 371234 336064 371240 336076
rect 371292 336064 371298 336116
rect 38746 335996 38752 336048
rect 38804 336036 38810 336048
rect 382366 336036 382372 336048
rect 38804 336008 382372 336036
rect 38804 335996 38810 336008
rect 382366 335996 382372 336008
rect 382424 335996 382430 336048
rect 82170 334568 82176 334620
rect 82228 334608 82234 334620
rect 178678 334608 178684 334620
rect 82228 334580 178684 334608
rect 82228 334568 82234 334580
rect 178678 334568 178684 334580
rect 178736 334568 178742 334620
rect 71314 331848 71320 331900
rect 71372 331888 71378 331900
rect 238754 331888 238760 331900
rect 71372 331860 238760 331888
rect 71372 331848 71378 331860
rect 238754 331848 238760 331860
rect 238812 331848 238818 331900
rect 68738 324300 68744 324352
rect 68796 324340 68802 324352
rect 579982 324340 579988 324352
rect 68796 324312 579988 324340
rect 68796 324300 68802 324312
rect 579982 324300 579988 324312
rect 580040 324300 580046 324352
rect 3418 318792 3424 318844
rect 3476 318832 3482 318844
rect 158714 318832 158720 318844
rect 3476 318804 158720 318832
rect 3476 318792 3482 318804
rect 158714 318792 158720 318804
rect 158772 318792 158778 318844
rect 70302 311856 70308 311908
rect 70360 311896 70366 311908
rect 580166 311896 580172 311908
rect 70360 311868 580172 311896
rect 70360 311856 70366 311868
rect 580166 311856 580172 311868
rect 580224 311856 580230 311908
rect 3418 304988 3424 305040
rect 3476 305028 3482 305040
rect 161474 305028 161480 305040
rect 3476 305000 161480 305028
rect 3476 304988 3482 305000
rect 161474 304988 161480 305000
rect 161532 304988 161538 305040
rect 67542 298120 67548 298172
rect 67600 298160 67606 298172
rect 580166 298160 580172 298172
rect 67600 298132 580172 298160
rect 67600 298120 67606 298132
rect 580166 298120 580172 298132
rect 580224 298120 580230 298172
rect 3418 292544 3424 292596
rect 3476 292584 3482 292596
rect 160094 292584 160100 292596
rect 3476 292556 160100 292584
rect 3476 292544 3482 292556
rect 160094 292544 160100 292556
rect 160152 292544 160158 292596
rect 66162 271872 66168 271924
rect 66220 271912 66226 271924
rect 580166 271912 580172 271924
rect 66220 271884 580172 271912
rect 66220 271872 66226 271884
rect 580166 271872 580172 271884
rect 580224 271872 580230 271924
rect 216582 269764 216588 269816
rect 216640 269804 216646 269816
rect 399570 269804 399576 269816
rect 216640 269776 399576 269804
rect 216640 269764 216646 269776
rect 399570 269764 399576 269776
rect 399628 269764 399634 269816
rect 10318 268404 10324 268456
rect 10376 268444 10382 268456
rect 139394 268444 139400 268456
rect 10376 268416 139400 268444
rect 10376 268404 10382 268416
rect 139394 268404 139400 268416
rect 139452 268404 139458 268456
rect 20070 268336 20076 268388
rect 20128 268376 20134 268388
rect 154574 268376 154580 268388
rect 20128 268348 154580 268376
rect 20128 268336 20134 268348
rect 154574 268336 154580 268348
rect 154632 268336 154638 268388
rect 108850 266976 108856 267028
rect 108908 267016 108914 267028
rect 215938 267016 215944 267028
rect 108908 266988 215944 267016
rect 108908 266976 108914 266988
rect 215938 266976 215944 266988
rect 215996 266976 216002 267028
rect 3050 266364 3056 266416
rect 3108 266404 3114 266416
rect 162854 266404 162860 266416
rect 3108 266376 162860 266404
rect 3108 266364 3114 266376
rect 162854 266364 162860 266376
rect 162912 266364 162918 266416
rect 32398 262896 32404 262948
rect 32456 262936 32462 262948
rect 149054 262936 149060 262948
rect 32456 262908 149060 262936
rect 32456 262896 32462 262908
rect 149054 262896 149060 262908
rect 149112 262896 149118 262948
rect 38838 262828 38844 262880
rect 38896 262868 38902 262880
rect 195974 262868 195980 262880
rect 38896 262840 195980 262868
rect 38896 262828 38902 262840
rect 195974 262828 195980 262840
rect 196032 262828 196038 262880
rect 66070 258068 66076 258120
rect 66128 258108 66134 258120
rect 580166 258108 580172 258120
rect 66128 258080 580172 258108
rect 66128 258068 66134 258080
rect 580166 258068 580172 258080
rect 580224 258068 580230 258120
rect 3418 253920 3424 253972
rect 3476 253960 3482 253972
rect 165614 253960 165620 253972
rect 3476 253932 165620 253960
rect 3476 253920 3482 253932
rect 165614 253920 165620 253932
rect 165672 253920 165678 253972
rect 86770 253172 86776 253224
rect 86828 253212 86834 253224
rect 231118 253212 231124 253224
rect 86828 253184 231124 253212
rect 86828 253172 86834 253184
rect 231118 253172 231124 253184
rect 231176 253172 231182 253224
rect 91002 252152 91008 252204
rect 91060 252192 91066 252204
rect 204990 252192 204996 252204
rect 91060 252164 204996 252192
rect 91060 252152 91066 252164
rect 204990 252152 204996 252164
rect 205048 252152 205054 252204
rect 106918 252084 106924 252136
rect 106976 252124 106982 252136
rect 229094 252124 229100 252136
rect 106976 252096 229100 252124
rect 106976 252084 106982 252096
rect 229094 252084 229100 252096
rect 229152 252084 229158 252136
rect 85482 252016 85488 252068
rect 85540 252056 85546 252068
rect 219434 252056 219440 252068
rect 85540 252028 219440 252056
rect 85540 252016 85546 252028
rect 219434 252016 219440 252028
rect 219492 252016 219498 252068
rect 79318 251948 79324 252000
rect 79376 251988 79382 252000
rect 213914 251988 213920 252000
rect 79376 251960 213920 251988
rect 79376 251948 79382 251960
rect 213914 251948 213920 251960
rect 213972 251948 213978 252000
rect 64782 251880 64788 251932
rect 64840 251920 64846 251932
rect 237926 251920 237932 251932
rect 64840 251892 237932 251920
rect 64840 251880 64846 251892
rect 237926 251880 237932 251892
rect 237984 251880 237990 251932
rect 35342 251812 35348 251864
rect 35400 251852 35406 251864
rect 393406 251852 393412 251864
rect 35400 251824 393412 251852
rect 35400 251812 35406 251824
rect 393406 251812 393412 251824
rect 393464 251812 393470 251864
rect 25498 250860 25504 250912
rect 25556 250900 25562 250912
rect 136634 250900 136640 250912
rect 25556 250872 136640 250900
rect 25556 250860 25562 250872
rect 136634 250860 136640 250872
rect 136692 250860 136698 250912
rect 119798 250792 119804 250844
rect 119856 250832 119862 250844
rect 282914 250832 282920 250844
rect 119856 250804 282920 250832
rect 119856 250792 119862 250804
rect 282914 250792 282920 250804
rect 282972 250792 282978 250844
rect 84286 250724 84292 250776
rect 84344 250764 84350 250776
rect 266998 250764 267004 250776
rect 84344 250736 267004 250764
rect 84344 250724 84350 250736
rect 266998 250724 267004 250736
rect 267056 250724 267062 250776
rect 35526 250656 35532 250708
rect 35584 250696 35590 250708
rect 369946 250696 369952 250708
rect 35584 250668 369952 250696
rect 35584 250656 35590 250668
rect 369946 250656 369952 250668
rect 370004 250656 370010 250708
rect 77294 250588 77300 250640
rect 77352 250628 77358 250640
rect 486418 250628 486424 250640
rect 77352 250600 486424 250628
rect 77352 250588 77358 250600
rect 486418 250588 486424 250600
rect 486476 250588 486482 250640
rect 71774 250520 71780 250572
rect 71832 250560 71838 250572
rect 483658 250560 483664 250572
rect 71832 250532 483664 250560
rect 71832 250520 71838 250532
rect 483658 250520 483664 250532
rect 483716 250520 483722 250572
rect 99374 250452 99380 250504
rect 99432 250492 99438 250504
rect 542354 250492 542360 250504
rect 99432 250464 542360 250492
rect 99432 250452 99438 250464
rect 542354 250452 542360 250464
rect 542412 250452 542418 250504
rect 117314 249704 117320 249756
rect 117372 249744 117378 249756
rect 201494 249744 201500 249756
rect 117372 249716 201500 249744
rect 117372 249704 117378 249716
rect 201494 249704 201500 249716
rect 201552 249704 201558 249756
rect 36630 249636 36636 249688
rect 36688 249676 36694 249688
rect 122834 249676 122840 249688
rect 36688 249648 122840 249676
rect 36688 249636 36694 249648
rect 122834 249636 122840 249648
rect 122892 249636 122898 249688
rect 100754 249568 100760 249620
rect 100812 249608 100818 249620
rect 189718 249608 189724 249620
rect 100812 249580 189724 249608
rect 100812 249568 100818 249580
rect 189718 249568 189724 249580
rect 189776 249568 189782 249620
rect 110414 249500 110420 249552
rect 110472 249540 110478 249552
rect 211798 249540 211804 249552
rect 110472 249512 211804 249540
rect 110472 249500 110478 249512
rect 211798 249500 211804 249512
rect 211856 249500 211862 249552
rect 95234 249432 95240 249484
rect 95292 249472 95298 249484
rect 196618 249472 196624 249484
rect 95292 249444 196624 249472
rect 95292 249432 95298 249444
rect 196618 249432 196624 249444
rect 196676 249432 196682 249484
rect 106274 249364 106280 249416
rect 106332 249404 106338 249416
rect 209038 249404 209044 249416
rect 106332 249376 209044 249404
rect 106332 249364 106338 249376
rect 209038 249364 209044 249376
rect 209096 249364 209102 249416
rect 102134 249296 102140 249348
rect 102192 249336 102198 249348
rect 204898 249336 204904 249348
rect 102192 249308 204904 249336
rect 102192 249296 102198 249308
rect 204898 249296 204904 249308
rect 204956 249296 204962 249348
rect 114554 249228 114560 249280
rect 114612 249268 114618 249280
rect 229738 249268 229744 249280
rect 114612 249240 229744 249268
rect 114612 249228 114618 249240
rect 229738 249228 229744 249240
rect 229796 249228 229802 249280
rect 86954 249160 86960 249212
rect 87012 249200 87018 249212
rect 226978 249200 226984 249212
rect 87012 249172 226984 249200
rect 87012 249160 87018 249172
rect 226978 249160 226984 249172
rect 227036 249160 227042 249212
rect 82814 249092 82820 249144
rect 82872 249132 82878 249144
rect 269758 249132 269764 249144
rect 82872 249104 269764 249132
rect 82872 249092 82878 249104
rect 269758 249092 269764 249104
rect 269816 249092 269822 249144
rect 35434 249024 35440 249076
rect 35492 249064 35498 249076
rect 380986 249064 380992 249076
rect 35492 249036 380992 249064
rect 35492 249024 35498 249036
rect 380986 249024 380992 249036
rect 381044 249024 381050 249076
rect 105722 248344 105728 248396
rect 105780 248384 105786 248396
rect 191098 248384 191104 248396
rect 105780 248356 191104 248384
rect 105780 248344 105786 248356
rect 191098 248344 191104 248356
rect 191156 248344 191162 248396
rect 98086 248276 98092 248328
rect 98144 248316 98150 248328
rect 185578 248316 185584 248328
rect 98144 248288 185584 248316
rect 98144 248276 98150 248288
rect 185578 248276 185584 248288
rect 185636 248276 185642 248328
rect 90358 248208 90364 248260
rect 90416 248248 90422 248260
rect 180058 248248 180064 248260
rect 90416 248220 180064 248248
rect 90416 248208 90422 248220
rect 180058 248208 180064 248220
rect 180116 248208 180122 248260
rect 91646 248140 91652 248192
rect 91704 248180 91710 248192
rect 200758 248180 200764 248192
rect 91704 248152 200764 248180
rect 91704 248140 91710 248152
rect 200758 248140 200764 248152
rect 200816 248140 200822 248192
rect 6178 248072 6184 248124
rect 6236 248112 6242 248124
rect 132586 248112 132592 248124
rect 6236 248084 132592 248112
rect 6236 248072 6242 248084
rect 132586 248072 132592 248084
rect 132644 248072 132650 248124
rect 86862 248004 86868 248056
rect 86920 248044 86926 248056
rect 241698 248044 241704 248056
rect 86920 248016 241704 248044
rect 86920 248004 86926 248016
rect 241698 248004 241704 248016
rect 241756 248004 241762 248056
rect 82630 247936 82636 247988
rect 82688 247976 82694 247988
rect 265618 247976 265624 247988
rect 82688 247948 265624 247976
rect 82688 247936 82694 247948
rect 265618 247936 265624 247948
rect 265676 247936 265682 247988
rect 80146 247868 80152 247920
rect 80204 247908 80210 247920
rect 268378 247908 268384 247920
rect 80204 247880 268384 247908
rect 80204 247868 80210 247880
rect 268378 247868 268384 247880
rect 268436 247868 268442 247920
rect 78858 247800 78864 247852
rect 78916 247840 78922 247852
rect 479518 247840 479524 247852
rect 78916 247812 479524 247840
rect 78916 247800 78922 247812
rect 479518 247800 479524 247812
rect 479576 247800 479582 247852
rect 75086 247732 75092 247784
rect 75144 247772 75150 247784
rect 482278 247772 482284 247784
rect 75144 247744 482284 247772
rect 75144 247732 75150 247744
rect 482278 247732 482284 247744
rect 482336 247732 482342 247784
rect 71222 247664 71228 247716
rect 71280 247704 71286 247716
rect 480898 247704 480904 247716
rect 71280 247676 480904 247704
rect 71280 247664 71286 247676
rect 480898 247664 480904 247676
rect 480956 247664 480962 247716
rect 109586 247596 109592 247648
rect 109644 247636 109650 247648
rect 193858 247636 193864 247648
rect 109644 247608 193864 247636
rect 109644 247596 109650 247608
rect 193858 247596 193864 247608
rect 193916 247596 193922 247648
rect 36814 247528 36820 247580
rect 36872 247568 36878 247580
rect 113174 247568 113180 247580
rect 36872 247540 113180 247568
rect 36872 247528 36878 247540
rect 113174 247528 113180 247540
rect 113232 247528 113238 247580
rect 94222 246848 94228 246900
rect 94280 246888 94286 246900
rect 182818 246888 182824 246900
rect 94280 246860 182824 246888
rect 94280 246848 94286 246860
rect 182818 246848 182824 246860
rect 182876 246848 182882 246900
rect 24762 246780 24768 246832
rect 24820 246820 24826 246832
rect 131298 246820 131304 246832
rect 24820 246792 131304 246820
rect 24820 246780 24826 246792
rect 131298 246780 131304 246792
rect 131356 246780 131362 246832
rect 93670 246712 93676 246764
rect 93728 246752 93734 246764
rect 208026 246752 208032 246764
rect 93728 246724 208032 246752
rect 93728 246712 93734 246724
rect 208026 246712 208032 246724
rect 208084 246712 208090 246764
rect 108942 246644 108948 246696
rect 109000 246684 109006 246696
rect 239306 246684 239312 246696
rect 109000 246656 239312 246684
rect 109000 246644 109006 246656
rect 239306 246644 239312 246656
rect 239364 246644 239370 246696
rect 60642 246576 60648 246628
rect 60700 246616 60706 246628
rect 192662 246616 192668 246628
rect 60700 246588 192668 246616
rect 60700 246576 60706 246588
rect 192662 246576 192668 246588
rect 192720 246576 192726 246628
rect 57882 246508 57888 246560
rect 57940 246548 57946 246560
rect 191374 246548 191380 246560
rect 57940 246520 191380 246548
rect 57940 246508 57946 246520
rect 191374 246508 191380 246520
rect 191432 246508 191438 246560
rect 38194 246440 38200 246492
rect 38252 246480 38258 246492
rect 186314 246480 186320 246492
rect 38252 246452 186320 246480
rect 38252 246440 38258 246452
rect 186314 246440 186320 246452
rect 186372 246440 186378 246492
rect 3694 246372 3700 246424
rect 3752 246412 3758 246424
rect 154298 246412 154304 246424
rect 3752 246384 154304 246412
rect 3752 246372 3758 246384
rect 154298 246372 154304 246384
rect 154356 246372 154362 246424
rect 38654 246304 38660 246356
rect 38712 246344 38718 246356
rect 199102 246344 199108 246356
rect 38712 246316 199108 246344
rect 38712 246304 38718 246316
rect 199102 246304 199108 246316
rect 199160 246304 199166 246356
rect 21358 245556 21364 245608
rect 21416 245596 21422 245608
rect 133874 245596 133880 245608
rect 21416 245568 133880 245596
rect 21416 245556 21422 245568
rect 133874 245556 133880 245568
rect 133932 245556 133938 245608
rect 31018 245488 31024 245540
rect 31076 245528 31082 245540
rect 145374 245528 145380 245540
rect 31076 245500 145380 245528
rect 31076 245488 31082 245500
rect 145374 245488 145380 245500
rect 145432 245488 145438 245540
rect 146202 245488 146208 245540
rect 146260 245528 146266 245540
rect 241606 245528 241612 245540
rect 146260 245500 241612 245528
rect 146260 245488 146266 245500
rect 241606 245488 241612 245500
rect 241664 245488 241670 245540
rect 33778 245420 33784 245472
rect 33836 245460 33842 245472
rect 153010 245460 153016 245472
rect 33836 245432 153016 245460
rect 33836 245420 33842 245432
rect 153010 245420 153016 245432
rect 153068 245420 153074 245472
rect 92934 245352 92940 245404
rect 92992 245392 92998 245404
rect 214558 245392 214564 245404
rect 92992 245364 214564 245392
rect 92992 245352 92998 245364
rect 214558 245352 214564 245364
rect 214616 245352 214622 245404
rect 102042 245284 102048 245336
rect 102100 245324 102106 245336
rect 239214 245324 239220 245336
rect 102100 245296 239220 245324
rect 102100 245284 102106 245296
rect 239214 245284 239220 245296
rect 239272 245284 239278 245336
rect 35250 245216 35256 245268
rect 35308 245256 35314 245268
rect 156874 245256 156880 245268
rect 35308 245228 156880 245256
rect 35308 245216 35314 245228
rect 156874 245216 156880 245228
rect 156932 245216 156938 245268
rect 205450 245216 205456 245268
rect 205508 245256 205514 245268
rect 349798 245256 349804 245268
rect 205508 245228 349804 245256
rect 205508 245216 205514 245228
rect 349798 245216 349804 245228
rect 349856 245216 349862 245268
rect 68830 245148 68836 245200
rect 68888 245188 68894 245200
rect 238938 245188 238944 245200
rect 68888 245160 238944 245188
rect 68888 245148 68894 245160
rect 238938 245148 238944 245160
rect 238996 245148 239002 245200
rect 8202 245080 8208 245132
rect 8260 245120 8266 245132
rect 130010 245120 130016 245132
rect 8260 245092 130016 245120
rect 8260 245080 8266 245092
rect 130010 245080 130016 245092
rect 130068 245080 130074 245132
rect 231026 245080 231032 245132
rect 231084 245120 231090 245132
rect 437474 245120 437480 245132
rect 231084 245092 437480 245120
rect 231084 245080 231090 245092
rect 437474 245080 437480 245092
rect 437532 245080 437538 245132
rect 39574 245012 39580 245064
rect 39632 245052 39638 245064
rect 89714 245052 89720 245064
rect 39632 245024 89720 245052
rect 39632 245012 39638 245024
rect 89714 245012 89720 245024
rect 89772 245012 89778 245064
rect 104434 245012 104440 245064
rect 104492 245052 104498 245064
rect 477494 245052 477500 245064
rect 104492 245024 477500 245052
rect 104492 245012 104498 245024
rect 477494 245012 477500 245024
rect 477552 245012 477558 245064
rect 73798 244944 73804 244996
rect 73856 244984 73862 244996
rect 485038 244984 485044 244996
rect 73856 244956 485044 244984
rect 73856 244944 73862 244956
rect 485038 244944 485044 244956
rect 485096 244944 485102 244996
rect 76374 244876 76380 244928
rect 76432 244916 76438 244928
rect 580442 244916 580448 244928
rect 76432 244888 580448 244916
rect 76432 244876 76438 244888
rect 580442 244876 580448 244888
rect 580500 244876 580506 244928
rect 28258 244808 28264 244860
rect 28316 244848 28322 244860
rect 141510 244848 141516 244860
rect 28316 244820 141516 244848
rect 28316 244808 28322 244820
rect 141510 244808 141516 244820
rect 141568 244808 141574 244860
rect 36906 244740 36912 244792
rect 36964 244780 36970 244792
rect 104894 244780 104900 244792
rect 36964 244752 104900 244780
rect 36964 244740 36970 244752
rect 104894 244740 104900 244752
rect 104952 244740 104958 244792
rect 112162 244740 112168 244792
rect 112220 244780 112226 244792
rect 220078 244780 220084 244792
rect 112220 244752 220084 244780
rect 112220 244740 112226 244752
rect 220078 244740 220084 244752
rect 220136 244740 220142 244792
rect 119982 244672 119988 244724
rect 120040 244712 120046 244724
rect 218054 244712 218060 244724
rect 120040 244684 218060 244712
rect 120040 244672 120046 244684
rect 218054 244672 218060 244684
rect 218112 244672 218118 244724
rect 117222 243924 117228 243976
rect 117280 243964 117286 243976
rect 197998 243964 198004 243976
rect 117280 243936 198004 243964
rect 117280 243924 117286 243936
rect 197998 243924 198004 243936
rect 198056 243924 198062 243976
rect 198090 243924 198096 243976
rect 198148 243964 198154 243976
rect 249058 243964 249064 243976
rect 198148 243936 249064 243964
rect 198148 243924 198154 243936
rect 249058 243924 249064 243936
rect 249116 243924 249122 243976
rect 15838 243856 15844 243908
rect 15896 243896 15902 243908
rect 136450 243896 136456 243908
rect 15896 243868 136456 243896
rect 15896 243856 15902 243868
rect 136450 243856 136456 243868
rect 136508 243856 136514 243908
rect 142062 243856 142068 243908
rect 142120 243896 142126 243908
rect 240594 243896 240600 243908
rect 142120 243868 240600 243896
rect 142120 243856 142126 243868
rect 240594 243856 240600 243868
rect 240652 243856 240658 243908
rect 13078 243788 13084 243840
rect 13136 243828 13142 243840
rect 144086 243828 144092 243840
rect 13136 243800 144092 243828
rect 13136 243788 13142 243800
rect 144086 243788 144092 243800
rect 144144 243788 144150 243840
rect 193950 243788 193956 243840
rect 194008 243828 194014 243840
rect 355318 243828 355324 243840
rect 194008 243800 355324 243828
rect 194008 243788 194014 243800
rect 355318 243788 355324 243800
rect 355376 243788 355382 243840
rect 113450 243720 113456 243772
rect 113508 243760 113514 243772
rect 299474 243760 299480 243772
rect 113508 243732 299480 243760
rect 113508 243720 113514 243732
rect 299474 243720 299480 243732
rect 299532 243720 299538 243772
rect 14458 243652 14464 243704
rect 14516 243692 14522 243704
rect 147950 243692 147956 243704
rect 14516 243664 147956 243692
rect 14516 243652 14522 243664
rect 147950 243652 147956 243664
rect 148008 243652 148014 243704
rect 225966 243652 225972 243704
rect 226024 243692 226030 243704
rect 430574 243692 430580 243704
rect 226024 243664 430580 243692
rect 226024 243652 226030 243664
rect 430574 243652 430580 243664
rect 430632 243652 430638 243704
rect 17218 243584 17224 243636
rect 17276 243624 17282 243636
rect 151814 243624 151820 243636
rect 17276 243596 151820 243624
rect 17276 243584 17282 243596
rect 151814 243584 151820 243596
rect 151872 243584 151878 243636
rect 236178 243584 236184 243636
rect 236236 243624 236242 243636
rect 445754 243624 445760 243636
rect 236236 243596 445760 243624
rect 236236 243584 236242 243596
rect 445754 243584 445760 243596
rect 445812 243584 445818 243636
rect 85482 243516 85488 243568
rect 85540 243556 85546 243568
rect 579614 243556 579620 243568
rect 85540 243528 579620 243556
rect 85540 243516 85546 243528
rect 579614 243516 579620 243528
rect 579672 243516 579678 243568
rect 15930 243448 15936 243500
rect 15988 243488 15994 243500
rect 167086 243488 167092 243500
rect 15988 243460 167092 243488
rect 15988 243448 15994 243460
rect 167086 243448 167092 243460
rect 167144 243448 167150 243500
rect 28258 243380 28264 243432
rect 28316 243420 28322 243432
rect 179874 243420 179880 243432
rect 28316 243392 179880 243420
rect 28316 243380 28322 243392
rect 179874 243380 179880 243392
rect 179932 243380 179938 243432
rect 17310 243312 17316 243364
rect 17368 243352 17374 243364
rect 170950 243352 170956 243364
rect 17368 243324 170956 243352
rect 17368 243312 17374 243324
rect 170950 243312 170956 243324
rect 171008 243312 171014 243364
rect 19978 243244 19984 243296
rect 20036 243284 20042 243296
rect 174814 243284 174820 243296
rect 20036 243256 174820 243284
rect 20036 243244 20042 243256
rect 174814 243244 174820 243256
rect 174872 243244 174878 243296
rect 21358 243176 21364 243228
rect 21416 243216 21422 243228
rect 182450 243216 182456 243228
rect 21416 243188 182456 243216
rect 21416 243176 21422 243188
rect 182450 243176 182456 243188
rect 182508 243176 182514 243228
rect 6178 243108 6184 243160
rect 6236 243148 6242 243160
rect 178586 243148 178592 243160
rect 6236 243120 178592 243148
rect 6236 243108 6242 243120
rect 178586 243108 178592 243120
rect 178644 243108 178650 243160
rect 48222 243040 48228 243092
rect 48280 243080 48286 243092
rect 268378 243080 268384 243092
rect 48280 243052 268384 243080
rect 48280 243040 48286 243052
rect 268378 243040 268384 243052
rect 268436 243040 268442 243092
rect 44358 242972 44364 243024
rect 44416 243012 44422 243024
rect 266998 243012 267004 243024
rect 44416 242984 267004 243012
rect 44416 242972 44422 242984
rect 266998 242972 267004 242984
rect 267056 242972 267062 243024
rect 41782 242904 41788 242956
rect 41840 242944 41846 242956
rect 273898 242944 273904 242956
rect 41840 242916 273904 242944
rect 41840 242904 41846 242916
rect 273898 242904 273904 242916
rect 273956 242904 273962 242956
rect 81434 242836 81440 242888
rect 81492 242876 81498 242888
rect 82722 242876 82728 242888
rect 81492 242848 82728 242876
rect 81492 242836 81498 242848
rect 82722 242836 82728 242848
rect 82780 242836 82786 242888
rect 82814 242836 82820 242888
rect 82872 242876 82878 242888
rect 84010 242876 84016 242888
rect 82872 242848 84016 242876
rect 82872 242836 82878 242848
rect 84010 242836 84016 242848
rect 84068 242836 84074 242888
rect 84286 242836 84292 242888
rect 84344 242876 84350 242888
rect 85298 242876 85304 242888
rect 84344 242848 85304 242876
rect 84344 242836 84350 242848
rect 85298 242836 85304 242848
rect 85356 242836 85362 242888
rect 86954 242836 86960 242888
rect 87012 242876 87018 242888
rect 87874 242876 87880 242888
rect 87012 242848 87880 242876
rect 87012 242836 87018 242848
rect 87874 242836 87880 242848
rect 87932 242836 87938 242888
rect 96798 242836 96804 242888
rect 96856 242876 96862 242888
rect 97902 242876 97908 242888
rect 96856 242848 97908 242876
rect 96856 242836 96862 242848
rect 97902 242836 97908 242848
rect 97960 242836 97966 242888
rect 99374 242836 99380 242888
rect 99432 242876 99438 242888
rect 100294 242876 100300 242888
rect 99432 242848 100300 242876
rect 99432 242836 99438 242848
rect 100294 242836 100300 242848
rect 100352 242836 100358 242888
rect 100754 242836 100760 242888
rect 100812 242876 100818 242888
rect 101950 242876 101956 242888
rect 100812 242848 101956 242876
rect 100812 242836 100818 242848
rect 101950 242836 101956 242848
rect 102008 242836 102014 242888
rect 102134 242836 102140 242888
rect 102192 242876 102198 242888
rect 103146 242876 103152 242888
rect 102192 242848 103152 242876
rect 102192 242836 102198 242848
rect 103146 242836 103152 242848
rect 103204 242836 103210 242888
rect 106274 242836 106280 242888
rect 106332 242876 106338 242888
rect 107010 242876 107016 242888
rect 106332 242848 107016 242876
rect 106332 242836 106338 242848
rect 107010 242836 107016 242848
rect 107068 242836 107074 242888
rect 117314 242836 117320 242888
rect 117372 242876 117378 242888
rect 118510 242876 118516 242888
rect 117372 242848 118516 242876
rect 117372 242836 117378 242848
rect 118510 242836 118516 242848
rect 118568 242836 118574 242888
rect 126238 242836 126244 242888
rect 126296 242876 126302 242888
rect 240502 242876 240508 242888
rect 126296 242848 240508 242876
rect 126296 242836 126302 242848
rect 240502 242836 240508 242848
rect 240560 242836 240566 242888
rect 79962 242768 79968 242820
rect 80020 242808 80026 242820
rect 80020 242780 233556 242808
rect 80020 242768 80026 242780
rect 96338 242700 96344 242752
rect 96396 242740 96402 242752
rect 232314 242740 232320 242752
rect 96396 242712 232320 242740
rect 96396 242700 96402 242712
rect 232314 242700 232320 242712
rect 232372 242700 232378 242752
rect 233528 242740 233556 242780
rect 233602 242768 233608 242820
rect 233660 242808 233666 242820
rect 234522 242808 234528 242820
rect 233660 242780 234528 242808
rect 233660 242768 233666 242780
rect 234522 242768 234528 242780
rect 234580 242768 234586 242820
rect 238110 242808 238116 242820
rect 234632 242780 238116 242808
rect 234632 242740 234660 242780
rect 238110 242768 238116 242780
rect 238168 242768 238174 242820
rect 233528 242712 234660 242740
rect 237466 242700 237472 242752
rect 237524 242740 237530 242752
rect 398098 242740 398104 242752
rect 237524 242712 398104 242740
rect 237524 242700 237530 242712
rect 398098 242700 398104 242712
rect 398156 242700 398162 242752
rect 99374 242632 99380 242684
rect 99432 242672 99438 242684
rect 100662 242672 100668 242684
rect 99432 242644 100668 242672
rect 99432 242632 99438 242644
rect 100662 242632 100668 242644
rect 100720 242632 100726 242684
rect 115934 242632 115940 242684
rect 115992 242672 115998 242684
rect 119798 242672 119804 242684
rect 115992 242644 119804 242672
rect 115992 242632 115998 242644
rect 119798 242632 119804 242644
rect 119856 242632 119862 242684
rect 177298 242632 177304 242684
rect 177356 242672 177362 242684
rect 215573 242675 215631 242681
rect 215573 242672 215585 242675
rect 177356 242644 215585 242672
rect 177356 242632 177362 242644
rect 215573 242641 215585 242644
rect 215619 242641 215631 242675
rect 215573 242635 215631 242641
rect 215662 242632 215668 242684
rect 215720 242672 215726 242684
rect 216582 242672 216588 242684
rect 215720 242644 216588 242672
rect 215720 242632 215726 242644
rect 216582 242632 216588 242644
rect 216640 242632 216646 242684
rect 220814 242632 220820 242684
rect 220872 242672 220878 242684
rect 220872 242644 224816 242672
rect 220872 242632 220878 242644
rect 175918 242564 175924 242616
rect 175976 242604 175982 242616
rect 224678 242604 224684 242616
rect 175976 242576 224684 242604
rect 175976 242564 175982 242576
rect 224678 242564 224684 242576
rect 224736 242564 224742 242616
rect 224788 242604 224816 242644
rect 225598 242632 225604 242684
rect 225656 242672 225662 242684
rect 227162 242672 227168 242684
rect 225656 242644 227168 242672
rect 225656 242632 225662 242644
rect 227162 242632 227168 242644
rect 227220 242632 227226 242684
rect 382918 242672 382924 242684
rect 227272 242644 382924 242672
rect 227272 242604 227300 242644
rect 382918 242632 382924 242644
rect 382976 242632 382982 242684
rect 224788 242576 227300 242604
rect 228450 242564 228456 242616
rect 228508 242604 228514 242616
rect 391198 242604 391204 242616
rect 228508 242576 391204 242604
rect 228508 242564 228514 242576
rect 391198 242564 391204 242576
rect 391256 242564 391262 242616
rect 64874 242496 64880 242548
rect 64932 242536 64938 242548
rect 66162 242536 66168 242548
rect 64932 242508 66168 242536
rect 64932 242496 64938 242508
rect 66162 242496 66168 242508
rect 66220 242496 66226 242548
rect 124950 242496 124956 242548
rect 125008 242536 125014 242548
rect 177022 242536 177028 242548
rect 125008 242508 177028 242536
rect 125008 242496 125014 242508
rect 177022 242496 177028 242508
rect 177080 242496 177086 242548
rect 204990 242496 204996 242548
rect 205048 242536 205054 242548
rect 206738 242536 206744 242548
rect 205048 242508 206744 242536
rect 205048 242496 205054 242508
rect 206738 242496 206744 242508
rect 206796 242496 206802 242548
rect 207658 242496 207664 242548
rect 207716 242536 207722 242548
rect 210602 242536 210608 242548
rect 207716 242508 210608 242536
rect 207716 242496 207722 242508
rect 210602 242496 210608 242508
rect 210660 242496 210666 242548
rect 211890 242496 211896 242548
rect 211948 242536 211954 242548
rect 375466 242536 375472 242548
rect 211948 242508 375472 242536
rect 211948 242496 211954 242508
rect 375466 242496 375472 242508
rect 375524 242496 375530 242548
rect 75178 242428 75184 242480
rect 75236 242468 75242 242480
rect 202874 242468 202880 242480
rect 75236 242440 202880 242468
rect 75236 242428 75242 242440
rect 202874 242428 202880 242440
rect 202932 242428 202938 242480
rect 209314 242428 209320 242480
rect 209372 242468 209378 242480
rect 373994 242468 374000 242480
rect 209372 242440 374000 242468
rect 209372 242428 209378 242440
rect 373994 242428 374000 242440
rect 374052 242428 374058 242480
rect 39758 242360 39764 242412
rect 39816 242400 39822 242412
rect 126238 242400 126244 242412
rect 39816 242372 126244 242400
rect 39816 242360 39822 242372
rect 126238 242360 126244 242372
rect 126296 242360 126302 242412
rect 200390 242360 200396 242412
rect 200448 242400 200454 242412
rect 366358 242400 366364 242412
rect 200448 242372 366364 242400
rect 200448 242360 200454 242372
rect 366358 242360 366364 242372
rect 366416 242360 366422 242412
rect 63586 242292 63592 242344
rect 63644 242332 63650 242344
rect 85482 242332 85488 242344
rect 63644 242304 85488 242332
rect 63644 242292 63650 242304
rect 85482 242292 85488 242304
rect 85540 242292 85546 242344
rect 123662 242292 123668 242344
rect 123720 242332 123726 242344
rect 176930 242332 176936 242344
rect 123720 242304 176936 242332
rect 123720 242292 123726 242304
rect 176930 242292 176936 242304
rect 176988 242292 176994 242344
rect 190086 242292 190092 242344
rect 190144 242332 190150 242344
rect 356054 242332 356060 242344
rect 190144 242304 356060 242332
rect 190144 242292 190150 242304
rect 356054 242292 356060 242304
rect 356112 242292 356118 242344
rect 36538 242224 36544 242276
rect 36596 242264 36602 242276
rect 125594 242264 125600 242276
rect 36596 242236 125600 242264
rect 36596 242224 36602 242236
rect 125594 242224 125600 242236
rect 125652 242224 125658 242276
rect 127434 242224 127440 242276
rect 127492 242264 127498 242276
rect 176654 242264 176660 242276
rect 127492 242236 176660 242264
rect 127492 242224 127498 242236
rect 176654 242224 176660 242236
rect 176712 242224 176718 242276
rect 188890 242224 188896 242276
rect 188948 242264 188954 242276
rect 363046 242264 363052 242276
rect 188948 242236 363052 242264
rect 188948 242224 188954 242236
rect 363046 242224 363052 242236
rect 363104 242224 363110 242276
rect 35250 242156 35256 242208
rect 35308 242196 35314 242208
rect 376754 242196 376760 242208
rect 35308 242168 376760 242196
rect 35308 242156 35314 242168
rect 376754 242156 376760 242168
rect 376812 242156 376818 242208
rect 133782 242088 133788 242140
rect 133840 242128 133846 242140
rect 239490 242128 239496 242140
rect 133840 242100 239496 242128
rect 133840 242088 133846 242100
rect 239490 242088 239496 242100
rect 239548 242088 239554 242140
rect 136542 242020 136548 242072
rect 136600 242060 136606 242072
rect 240134 242060 240140 242072
rect 136600 242032 240140 242060
rect 136600 242020 136606 242032
rect 240134 242020 240140 242032
rect 240192 242020 240198 242072
rect 61010 241952 61016 242004
rect 61068 241992 61074 242004
rect 96522 241992 96528 242004
rect 61068 241964 96528 241992
rect 61068 241952 61074 241964
rect 96522 241952 96528 241964
rect 96580 241952 96586 242004
rect 178678 241952 178684 242004
rect 178736 241992 178742 242004
rect 218238 241992 218244 242004
rect 178736 241964 218244 241992
rect 178736 241952 178742 241964
rect 218238 241952 218244 241964
rect 218296 241952 218302 242004
rect 234890 241952 234896 242004
rect 234948 241992 234954 242004
rect 247678 241992 247684 242004
rect 234948 241964 247684 241992
rect 234948 241952 234954 241964
rect 247678 241952 247684 241964
rect 247736 241952 247742 242004
rect 53282 241884 53288 241936
rect 53340 241924 53346 241936
rect 128814 241924 128820 241936
rect 53340 241896 128820 241924
rect 53340 241884 53346 241896
rect 128814 241884 128820 241896
rect 128872 241884 128878 241936
rect 173158 241884 173164 241936
rect 173216 241924 173222 241936
rect 201586 241924 201592 241936
rect 173216 241896 201592 241924
rect 173216 241884 173222 241896
rect 201586 241884 201592 241896
rect 201644 241884 201650 241936
rect 215573 241927 215631 241933
rect 215573 241893 215585 241927
rect 215619 241924 215631 241927
rect 216950 241924 216956 241936
rect 215619 241896 216956 241924
rect 215619 241893 215631 241896
rect 215573 241887 215631 241893
rect 216950 241884 216956 241896
rect 217008 241884 217014 241936
rect 62298 241816 62304 241868
rect 62356 241856 62362 241868
rect 178034 241856 178040 241868
rect 62356 241828 178040 241856
rect 62356 241816 62362 241828
rect 178034 241816 178040 241828
rect 178092 241816 178098 241868
rect 58434 241748 58440 241800
rect 58492 241788 58498 241800
rect 177390 241788 177396 241800
rect 58492 241760 177396 241788
rect 58492 241748 58498 241760
rect 177390 241748 177396 241760
rect 177448 241748 177454 241800
rect 46934 241680 46940 241732
rect 46992 241720 46998 241732
rect 175182 241720 175188 241732
rect 46992 241692 175188 241720
rect 46992 241680 46998 241692
rect 175182 241680 175188 241692
rect 175240 241680 175246 241732
rect 3418 241612 3424 241664
rect 3476 241652 3482 241664
rect 164510 241652 164516 241664
rect 3476 241624 164516 241652
rect 3476 241612 3482 241624
rect 164510 241612 164516 241624
rect 164568 241612 164574 241664
rect 13078 241544 13084 241596
rect 13136 241584 13142 241596
rect 181162 241584 181168 241596
rect 13136 241556 181168 241584
rect 13136 241544 13142 241556
rect 181162 241544 181168 241556
rect 181220 241544 181226 241596
rect 14458 241476 14464 241528
rect 14516 241516 14522 241528
rect 185026 241516 185032 241528
rect 14516 241488 185032 241516
rect 14516 241476 14522 241488
rect 185026 241476 185032 241488
rect 185084 241476 185090 241528
rect 38562 241408 38568 241460
rect 38620 241448 38626 241460
rect 39298 241448 39304 241460
rect 38620 241420 39304 241448
rect 38620 241408 38626 241420
rect 39298 241408 39304 241420
rect 39356 241408 39362 241460
rect 39390 241408 39396 241460
rect 39448 241448 39454 241460
rect 74626 241448 74632 241460
rect 39448 241420 74632 241448
rect 39448 241408 39454 241420
rect 74626 241408 74632 241420
rect 74684 241408 74690 241460
rect 39114 241340 39120 241392
rect 39172 241380 39178 241392
rect 85666 241380 85672 241392
rect 39172 241352 85672 241380
rect 39172 241340 39178 241352
rect 85666 241340 85672 241352
rect 85724 241340 85730 241392
rect 39206 241272 39212 241324
rect 39264 241312 39270 241324
rect 87046 241312 87052 241324
rect 39264 241284 87052 241312
rect 39264 241272 39270 241284
rect 87046 241272 87052 241284
rect 87104 241272 87110 241324
rect 99098 241272 99104 241324
rect 99156 241312 99162 241324
rect 238846 241312 238852 241324
rect 99156 241284 238852 241312
rect 99156 241272 99162 241284
rect 238846 241272 238852 241284
rect 238904 241272 238910 241324
rect 39482 241204 39488 241256
rect 39540 241244 39546 241256
rect 91186 241244 91192 241256
rect 39540 241216 91192 241244
rect 39540 241204 39546 241216
rect 91186 241204 91192 241216
rect 91244 241204 91250 241256
rect 92382 241204 92388 241256
rect 92440 241244 92446 241256
rect 238018 241244 238024 241256
rect 92440 241216 238024 241244
rect 92440 241204 92446 241216
rect 238018 241204 238024 241216
rect 238076 241204 238082 241256
rect 68922 241136 68928 241188
rect 68980 241176 68986 241188
rect 239122 241176 239128 241188
rect 68980 241148 239128 241176
rect 68980 241136 68986 241148
rect 239122 241136 239128 241148
rect 239180 241136 239186 241188
rect 38838 241068 38844 241120
rect 38896 241108 38902 241120
rect 365714 241108 365720 241120
rect 38896 241080 365720 241108
rect 38896 241068 38902 241080
rect 365714 241068 365720 241080
rect 365772 241068 365778 241120
rect 36998 241000 37004 241052
rect 37056 241040 37062 241052
rect 367186 241040 367192 241052
rect 37056 241012 367192 241040
rect 37056 241000 37062 241012
rect 367186 241000 367192 241012
rect 367244 241000 367250 241052
rect 38102 240932 38108 240984
rect 38160 240972 38166 240984
rect 368474 240972 368480 240984
rect 38160 240944 368480 240972
rect 38160 240932 38166 240944
rect 368474 240932 368480 240944
rect 368532 240932 368538 240984
rect 37734 240864 37740 240916
rect 37792 240904 37798 240916
rect 381538 240904 381544 240916
rect 37792 240876 381544 240904
rect 37792 240864 37798 240876
rect 381538 240864 381544 240876
rect 381596 240864 381602 240916
rect 36722 240796 36728 240848
rect 36780 240836 36786 240848
rect 412634 240836 412640 240848
rect 36780 240808 412640 240836
rect 36780 240796 36786 240808
rect 412634 240796 412640 240808
rect 412692 240796 412698 240848
rect 61378 240728 61384 240780
rect 61436 240768 61442 240780
rect 240410 240768 240416 240780
rect 61436 240740 240416 240768
rect 61436 240728 61442 240740
rect 240410 240728 240416 240740
rect 240468 240728 240474 240780
rect 39022 240116 39028 240168
rect 39080 240156 39086 240168
rect 39390 240156 39396 240168
rect 39080 240128 39396 240156
rect 39080 240116 39086 240128
rect 39390 240116 39396 240128
rect 39448 240116 39454 240168
rect 168466 240048 168472 240100
rect 168524 240088 168530 240100
rect 580166 240088 580172 240100
rect 168524 240060 580172 240088
rect 168524 240048 168530 240060
rect 580166 240048 580172 240060
rect 580224 240048 580230 240100
rect 38010 239980 38016 240032
rect 38068 240020 38074 240032
rect 42058 240020 42064 240032
rect 38068 239992 42064 240020
rect 38068 239980 38074 239992
rect 42058 239980 42064 239992
rect 42116 239980 42122 240032
rect 236638 239980 236644 240032
rect 236696 240020 236702 240032
rect 237834 240020 237840 240032
rect 236696 239992 237840 240020
rect 236696 239980 236702 239992
rect 237834 239980 237840 239992
rect 237892 239980 237898 240032
rect 237929 240023 237987 240029
rect 237929 239989 237941 240023
rect 237975 240020 237987 240023
rect 240870 240020 240876 240032
rect 237975 239992 240876 240020
rect 237975 239989 237987 239992
rect 237929 239983 237987 239989
rect 240870 239980 240876 239992
rect 240928 239980 240934 240032
rect 37918 239912 37924 239964
rect 37976 239952 37982 239964
rect 46198 239952 46204 239964
rect 37976 239924 46204 239952
rect 37976 239912 37982 239924
rect 46198 239912 46204 239924
rect 46256 239912 46262 239964
rect 48869 239955 48927 239961
rect 48869 239921 48881 239955
rect 48915 239952 48927 239955
rect 171870 239952 171876 239964
rect 48915 239924 55214 239952
rect 171831 239924 171876 239952
rect 48915 239921 48927 239924
rect 48869 239915 48927 239921
rect 37826 239844 37832 239896
rect 37884 239884 37890 239896
rect 48958 239884 48964 239896
rect 37884 239856 48964 239884
rect 37884 239844 37890 239856
rect 48958 239844 48964 239856
rect 49016 239844 49022 239896
rect 50338 239884 50344 239896
rect 49068 239856 50344 239884
rect 33778 239776 33784 239828
rect 33836 239816 33842 239828
rect 48869 239819 48927 239825
rect 48869 239816 48881 239819
rect 33836 239788 48881 239816
rect 33836 239776 33842 239788
rect 48869 239785 48881 239788
rect 48915 239785 48927 239819
rect 48869 239779 48927 239785
rect 39390 239708 39396 239760
rect 39448 239748 39454 239760
rect 39574 239748 39580 239760
rect 39448 239720 39580 239748
rect 39448 239708 39454 239720
rect 39574 239708 39580 239720
rect 39632 239708 39638 239760
rect 40126 239708 40132 239760
rect 40184 239748 40190 239760
rect 43438 239748 43444 239760
rect 40184 239720 43444 239748
rect 40184 239708 40190 239720
rect 43438 239708 43444 239720
rect 43496 239708 43502 239760
rect 43533 239751 43591 239757
rect 43533 239717 43545 239751
rect 43579 239748 43591 239751
rect 49068 239748 49096 239856
rect 50338 239844 50344 239856
rect 50396 239844 50402 239896
rect 55186 239816 55214 239924
rect 171870 239912 171876 239924
rect 171928 239912 171934 239964
rect 236730 239912 236736 239964
rect 236788 239952 236794 239964
rect 240318 239952 240324 239964
rect 236788 239924 240324 239952
rect 236788 239912 236794 239924
rect 240318 239912 240324 239924
rect 240376 239912 240382 239964
rect 139302 239844 139308 239896
rect 139360 239884 139366 239896
rect 239030 239884 239036 239896
rect 139360 239856 239036 239884
rect 139360 239844 139366 239856
rect 239030 239844 239036 239856
rect 239088 239844 239094 239896
rect 183554 239816 183560 239828
rect 55186 239788 183560 239816
rect 183554 239776 183560 239788
rect 183612 239776 183618 239828
rect 232498 239776 232504 239828
rect 232556 239816 232562 239828
rect 237929 239819 237987 239825
rect 237929 239816 237941 239819
rect 232556 239788 237941 239816
rect 232556 239776 232562 239788
rect 237929 239785 237941 239788
rect 237975 239785 237987 239819
rect 237929 239779 237987 239785
rect 49602 239748 49608 239760
rect 43579 239720 49096 239748
rect 49563 239720 49608 239748
rect 43579 239717 43591 239720
rect 43533 239711 43591 239717
rect 49602 239708 49608 239720
rect 49660 239708 49666 239760
rect 52362 239748 52368 239760
rect 52323 239720 52368 239748
rect 52362 239708 52368 239720
rect 52420 239708 52426 239760
rect 54846 239748 54852 239760
rect 54807 239720 54852 239748
rect 54846 239708 54852 239720
rect 54904 239708 54910 239760
rect 56226 239748 56232 239760
rect 56187 239720 56232 239748
rect 56226 239708 56232 239720
rect 56284 239708 56290 239760
rect 57514 239748 57520 239760
rect 57475 239720 57520 239748
rect 57514 239708 57520 239720
rect 57572 239708 57578 239760
rect 57698 239748 57704 239760
rect 57659 239720 57704 239748
rect 57698 239708 57704 239720
rect 57756 239708 57762 239760
rect 59170 239748 59176 239760
rect 59131 239720 59176 239748
rect 59170 239708 59176 239720
rect 59228 239708 59234 239760
rect 60090 239748 60096 239760
rect 60051 239720 60096 239748
rect 60090 239708 60096 239720
rect 60148 239708 60154 239760
rect 62114 239748 62120 239760
rect 62075 239720 62120 239748
rect 62114 239708 62120 239720
rect 62172 239708 62178 239760
rect 73430 239748 73436 239760
rect 73391 239720 73436 239748
rect 73430 239708 73436 239720
rect 73488 239708 73494 239760
rect 75822 239748 75828 239760
rect 75783 239720 75828 239748
rect 75822 239708 75828 239720
rect 75880 239708 75886 239760
rect 82906 239748 82912 239760
rect 82867 239720 82912 239748
rect 82906 239708 82912 239720
rect 82964 239708 82970 239760
rect 96522 239708 96528 239760
rect 96580 239748 96586 239760
rect 97445 239751 97503 239757
rect 97445 239748 97457 239751
rect 96580 239720 97457 239748
rect 96580 239708 96586 239720
rect 97445 239717 97457 239720
rect 97491 239717 97503 239751
rect 128814 239748 128820 239760
rect 128775 239720 128820 239748
rect 97445 239711 97503 239717
rect 128814 239708 128820 239720
rect 128872 239708 128878 239760
rect 173158 239748 173164 239760
rect 161446 239720 173164 239748
rect 31018 239640 31024 239692
rect 31076 239680 31082 239692
rect 161446 239680 161474 239720
rect 173158 239708 173164 239720
rect 173216 239708 173222 239760
rect 175182 239708 175188 239760
rect 175240 239748 175246 239760
rect 175240 239720 175964 239748
rect 175240 239708 175246 239720
rect 168466 239680 168472 239692
rect 31076 239652 161474 239680
rect 168427 239652 168472 239680
rect 31076 239640 31082 239652
rect 168466 239640 168472 239652
rect 168524 239640 168530 239692
rect 169294 239680 169300 239692
rect 169255 239652 169300 239680
rect 169294 239640 169300 239652
rect 169352 239640 169358 239692
rect 175734 239680 175740 239692
rect 171106 239652 175740 239680
rect 25498 239572 25504 239624
rect 25556 239612 25562 239624
rect 171106 239612 171134 239652
rect 175734 239640 175740 239652
rect 175792 239640 175798 239692
rect 25556 239584 171134 239612
rect 175936 239612 175964 239720
rect 178034 239708 178040 239760
rect 178092 239748 178098 239760
rect 580626 239748 580632 239760
rect 178092 239720 580632 239748
rect 178092 239708 178098 239720
rect 580626 239708 580632 239720
rect 580684 239708 580690 239760
rect 177022 239680 177028 239692
rect 176983 239652 177028 239680
rect 177022 239640 177028 239652
rect 177080 239640 177086 239692
rect 177390 239640 177396 239692
rect 177448 239680 177454 239692
rect 580534 239680 580540 239692
rect 177448 239652 580540 239680
rect 177448 239640 177454 239652
rect 580534 239640 580540 239652
rect 580592 239640 580598 239692
rect 175936 239584 180794 239612
rect 25556 239572 25562 239584
rect 24118 239504 24124 239556
rect 24176 239544 24182 239556
rect 171873 239547 171931 239553
rect 171873 239544 171885 239547
rect 24176 239516 171885 239544
rect 24176 239504 24182 239516
rect 171873 239513 171885 239516
rect 171919 239513 171931 239547
rect 180766 239544 180794 239584
rect 580258 239544 580264 239556
rect 180766 239516 580264 239544
rect 171873 239507 171931 239513
rect 580258 239504 580264 239516
rect 580316 239504 580322 239556
rect 40218 239436 40224 239488
rect 40276 239476 40282 239488
rect 43533 239479 43591 239485
rect 43533 239476 43545 239479
rect 40276 239448 43545 239476
rect 40276 239436 40282 239448
rect 43533 239445 43545 239448
rect 43579 239445 43591 239479
rect 43533 239439 43591 239445
rect 43625 239479 43683 239485
rect 43625 239445 43637 239479
rect 43671 239476 43683 239479
rect 62117 239479 62175 239485
rect 62117 239476 62129 239479
rect 43671 239448 62129 239476
rect 43671 239445 43683 239448
rect 43625 239439 43683 239445
rect 62117 239445 62129 239448
rect 62163 239445 62175 239479
rect 62117 239439 62175 239445
rect 128817 239479 128875 239485
rect 128817 239445 128829 239479
rect 128863 239476 128875 239479
rect 580442 239476 580448 239488
rect 128863 239448 580448 239476
rect 128863 239445 128875 239448
rect 128817 239439 128875 239445
rect 580442 239436 580448 239448
rect 580500 239436 580506 239488
rect 38930 239368 38936 239420
rect 38988 239408 38994 239420
rect 82909 239411 82967 239417
rect 82909 239408 82921 239411
rect 38988 239380 82921 239408
rect 38988 239368 38994 239380
rect 82909 239377 82921 239380
rect 82955 239377 82967 239411
rect 82909 239371 82967 239377
rect 97445 239411 97503 239417
rect 97445 239377 97457 239411
rect 97491 239408 97503 239411
rect 580350 239408 580356 239420
rect 97491 239380 580356 239408
rect 97491 239377 97503 239380
rect 97445 239371 97503 239377
rect 580350 239368 580356 239380
rect 580408 239368 580414 239420
rect 10318 239300 10324 239352
rect 10376 239340 10382 239352
rect 169297 239343 169355 239349
rect 169297 239340 169309 239343
rect 10376 239312 169309 239340
rect 10376 239300 10382 239312
rect 169297 239309 169309 239312
rect 169343 239309 169355 239343
rect 169297 239303 169355 239309
rect 7558 239232 7564 239284
rect 7616 239272 7622 239284
rect 168469 239275 168527 239281
rect 168469 239272 168481 239275
rect 7616 239244 168481 239272
rect 7616 239232 7622 239244
rect 168469 239241 168481 239244
rect 168515 239241 168527 239275
rect 168469 239235 168527 239241
rect 3418 239164 3424 239216
rect 3476 239204 3482 239216
rect 177025 239207 177083 239213
rect 177025 239204 177037 239207
rect 3476 239176 177037 239204
rect 3476 239164 3482 239176
rect 177025 239173 177037 239176
rect 177071 239173 177083 239207
rect 177025 239167 177083 239173
rect 38654 239096 38660 239148
rect 38712 239136 38718 239148
rect 43625 239139 43683 239145
rect 43625 239136 43637 239139
rect 38712 239108 43637 239136
rect 38712 239096 38718 239108
rect 43625 239105 43637 239108
rect 43671 239105 43683 239139
rect 43625 239099 43683 239105
rect 60093 239139 60151 239145
rect 60093 239105 60105 239139
rect 60139 239136 60151 239139
rect 272518 239136 272524 239148
rect 60139 239108 272524 239136
rect 60139 239105 60151 239108
rect 60093 239099 60151 239105
rect 272518 239096 272524 239108
rect 272576 239096 272582 239148
rect 56229 239071 56287 239077
rect 56229 239037 56241 239071
rect 56275 239068 56287 239071
rect 269758 239068 269764 239080
rect 56275 239040 269764 239068
rect 56275 239037 56287 239040
rect 56229 239031 56287 239037
rect 269758 239028 269764 239040
rect 269816 239028 269822 239080
rect 57517 239003 57575 239009
rect 57517 238969 57529 239003
rect 57563 239000 57575 239003
rect 280798 239000 280804 239012
rect 57563 238972 280804 239000
rect 57563 238969 57575 238972
rect 57517 238963 57575 238969
rect 280798 238960 280804 238972
rect 280856 238960 280862 239012
rect 49605 238935 49663 238941
rect 49605 238901 49617 238935
rect 49651 238932 49663 238935
rect 279418 238932 279424 238944
rect 49651 238904 279424 238932
rect 49651 238901 49663 238904
rect 49605 238895 49663 238901
rect 279418 238892 279424 238904
rect 279476 238892 279482 238944
rect 54849 238867 54907 238873
rect 54849 238833 54861 238867
rect 54895 238864 54907 238867
rect 284938 238864 284944 238876
rect 54895 238836 284944 238864
rect 54895 238833 54907 238836
rect 54849 238827 54907 238833
rect 284938 238824 284944 238836
rect 284996 238824 285002 238876
rect 52365 238799 52423 238805
rect 52365 238765 52377 238799
rect 52411 238796 52423 238799
rect 341518 238796 341524 238808
rect 52411 238768 341524 238796
rect 52411 238765 52423 238768
rect 52365 238759 52423 238765
rect 341518 238756 341524 238768
rect 341576 238756 341582 238808
rect 38562 238688 38568 238740
rect 38620 238728 38626 238740
rect 40218 238728 40224 238740
rect 38620 238700 40224 238728
rect 38620 238688 38626 238700
rect 40218 238688 40224 238700
rect 40276 238688 40282 238740
rect 241146 238688 241152 238740
rect 241204 238728 241210 238740
rect 364978 238728 364984 238740
rect 241204 238700 364984 238728
rect 241204 238688 241210 238700
rect 364978 238688 364984 238700
rect 365036 238688 365042 238740
rect 59173 238323 59231 238329
rect 59173 238289 59185 238323
rect 59219 238320 59231 238323
rect 73433 238323 73491 238329
rect 73433 238320 73445 238323
rect 59219 238292 73445 238320
rect 59219 238289 59231 238292
rect 59173 238283 59231 238289
rect 73433 238289 73445 238292
rect 73479 238289 73491 238323
rect 73433 238283 73491 238289
rect 57701 238255 57759 238261
rect 57701 238221 57713 238255
rect 57747 238252 57759 238255
rect 75825 238255 75883 238261
rect 75825 238252 75837 238255
rect 57747 238224 75837 238252
rect 57747 238221 57759 238224
rect 57701 238215 57759 238221
rect 75825 238221 75837 238224
rect 75871 238221 75883 238255
rect 75825 238215 75883 238221
rect 38286 238144 38292 238196
rect 38344 238184 38350 238196
rect 357434 238184 357440 238196
rect 38344 238156 357440 238184
rect 38344 238144 38350 238156
rect 357434 238144 357440 238156
rect 357492 238144 357498 238196
rect 580350 235492 580356 235544
rect 580408 235532 580414 235544
rect 580718 235532 580724 235544
rect 580408 235504 580724 235532
rect 580408 235492 580414 235504
rect 580718 235492 580724 235504
rect 580776 235492 580782 235544
rect 38194 232772 38200 232824
rect 38252 232812 38258 232824
rect 40402 232812 40408 232824
rect 38252 232784 40408 232812
rect 38252 232772 38258 232784
rect 40402 232772 40408 232784
rect 40460 232772 40466 232824
rect 38286 231956 38292 232008
rect 38344 231996 38350 232008
rect 38562 231996 38568 232008
rect 38344 231968 38568 231996
rect 38344 231956 38350 231968
rect 38562 231956 38568 231968
rect 38620 231956 38626 232008
rect 238294 229032 238300 229084
rect 238352 229072 238358 229084
rect 240594 229072 240600 229084
rect 238352 229044 240600 229072
rect 238352 229032 238358 229044
rect 240594 229032 240600 229044
rect 240652 229032 240658 229084
rect 240226 226992 240232 227044
rect 240284 227032 240290 227044
rect 240410 227032 240416 227044
rect 240284 227004 240416 227032
rect 240284 226992 240290 227004
rect 240410 226992 240416 227004
rect 240468 226992 240474 227044
rect 240318 226040 240324 226092
rect 240376 226040 240382 226092
rect 240336 225888 240364 226040
rect 240318 225836 240324 225888
rect 240376 225836 240382 225888
rect 239398 224748 239404 224800
rect 239456 224788 239462 224800
rect 240410 224788 240416 224800
rect 239456 224760 240416 224788
rect 239456 224748 239462 224760
rect 240410 224748 240416 224760
rect 240468 224748 240474 224800
rect 3326 215228 3332 215280
rect 3384 215268 3390 215280
rect 15930 215268 15936 215280
rect 3384 215240 15936 215268
rect 3384 215228 3390 215240
rect 15930 215228 15936 215240
rect 15988 215228 15994 215280
rect 241238 213868 241244 213920
rect 241296 213908 241302 213920
rect 251818 213908 251824 213920
rect 241296 213880 251824 213908
rect 241296 213868 241302 213880
rect 251818 213868 251824 213880
rect 251876 213868 251882 213920
rect 241422 208292 241428 208344
rect 241480 208332 241486 208344
rect 388438 208332 388444 208344
rect 241480 208304 388444 208332
rect 241480 208292 241486 208304
rect 388438 208292 388444 208304
rect 388496 208292 388502 208344
rect 272518 206932 272524 206984
rect 272576 206972 272582 206984
rect 579798 206972 579804 206984
rect 272576 206944 579804 206972
rect 272576 206932 272582 206944
rect 579798 206932 579804 206944
rect 579856 206932 579862 206984
rect 285674 204892 285680 204944
rect 285732 204932 285738 204944
rect 427814 204932 427820 204944
rect 285732 204904 427820 204932
rect 285732 204892 285738 204904
rect 427814 204892 427820 204904
rect 427872 204892 427878 204944
rect 3050 202784 3056 202836
rect 3108 202824 3114 202836
rect 10318 202824 10324 202836
rect 3108 202796 10324 202824
rect 3108 202784 3114 202796
rect 10318 202784 10324 202796
rect 10376 202784 10382 202836
rect 241422 202784 241428 202836
rect 241480 202824 241486 202836
rect 285674 202824 285680 202836
rect 241480 202796 285680 202824
rect 241480 202784 241486 202796
rect 285674 202784 285680 202796
rect 285732 202784 285738 202836
rect 241422 198636 241428 198688
rect 241480 198676 241486 198688
rect 387058 198676 387064 198688
rect 241480 198648 387064 198676
rect 241480 198636 241486 198648
rect 387058 198636 387064 198648
rect 387116 198636 387122 198688
rect 238202 195916 238208 195968
rect 238260 195956 238266 195968
rect 240134 195956 240140 195968
rect 238260 195928 240140 195956
rect 238260 195916 238266 195928
rect 240134 195916 240140 195928
rect 240192 195916 240198 195968
rect 280798 193128 280804 193180
rect 280856 193168 280862 193180
rect 579614 193168 579620 193180
rect 280856 193140 579620 193168
rect 280856 193128 280862 193140
rect 579614 193128 579620 193140
rect 579672 193128 579678 193180
rect 3510 188844 3516 188896
rect 3568 188884 3574 188896
rect 7558 188884 7564 188896
rect 3568 188856 7564 188884
rect 3568 188844 3574 188856
rect 7558 188844 7564 188856
rect 7616 188844 7622 188896
rect 241422 187620 241428 187672
rect 241480 187660 241486 187672
rect 417418 187660 417424 187672
rect 241480 187632 417424 187660
rect 241480 187620 241486 187632
rect 417418 187620 417424 187632
rect 417476 187620 417482 187672
rect 285674 185580 285680 185632
rect 285732 185620 285738 185632
rect 415394 185620 415400 185632
rect 285732 185592 415400 185620
rect 285732 185580 285738 185592
rect 415394 185580 415400 185592
rect 415452 185580 415458 185632
rect 241422 183472 241428 183524
rect 241480 183512 241486 183524
rect 285674 183512 285680 183524
rect 241480 183484 285680 183512
rect 241480 183472 241486 183484
rect 285674 183472 285680 183484
rect 285732 183472 285738 183524
rect 241238 173612 241244 173664
rect 241296 173652 241302 173664
rect 244918 173652 244924 173664
rect 241296 173624 244924 173652
rect 241296 173612 241302 173624
rect 244918 173612 244924 173624
rect 244976 173612 244982 173664
rect 35618 169464 35624 169516
rect 35676 169504 35682 169516
rect 37826 169504 37832 169516
rect 35676 169476 37832 169504
rect 35676 169464 35682 169476
rect 37826 169464 37832 169476
rect 37884 169464 37890 169516
rect 269758 166948 269764 167000
rect 269816 166988 269822 167000
rect 580166 166988 580172 167000
rect 269816 166960 580172 166988
rect 269816 166948 269822 166960
rect 580166 166948 580172 166960
rect 580224 166948 580230 167000
rect 3234 164160 3240 164212
rect 3292 164200 3298 164212
rect 17310 164200 17316 164212
rect 3292 164172 17316 164200
rect 3292 164160 3298 164172
rect 17310 164160 17316 164172
rect 17368 164160 17374 164212
rect 241054 158040 241060 158092
rect 241112 158080 241118 158092
rect 243538 158080 243544 158092
rect 241112 158052 243544 158080
rect 241112 158040 241118 158052
rect 243538 158040 243544 158052
rect 243596 158040 243602 158092
rect 35250 151716 35256 151768
rect 35308 151756 35314 151768
rect 37734 151756 37740 151768
rect 35308 151728 37740 151756
rect 35308 151716 35314 151728
rect 37734 151716 37740 151728
rect 37792 151716 37798 151768
rect 3510 150356 3516 150408
rect 3568 150396 3574 150408
rect 31018 150396 31024 150408
rect 3568 150368 31024 150396
rect 3568 150356 3574 150368
rect 31018 150356 31024 150368
rect 31076 150356 31082 150408
rect 241146 143488 241152 143540
rect 241204 143528 241210 143540
rect 371878 143528 371884 143540
rect 241204 143500 371884 143528
rect 241204 143488 241210 143500
rect 371878 143488 371884 143500
rect 371936 143488 371942 143540
rect 284938 139340 284944 139392
rect 284996 139380 285002 139392
rect 580166 139380 580172 139392
rect 284996 139352 580172 139380
rect 284996 139340 285002 139352
rect 580166 139340 580172 139352
rect 580224 139340 580230 139392
rect 3510 137912 3516 137964
rect 3568 137952 3574 137964
rect 24118 137952 24124 137964
rect 3568 137924 24124 137952
rect 3568 137912 3574 137924
rect 24118 137912 24124 137924
rect 24176 137912 24182 137964
rect 241422 137912 241428 137964
rect 241480 137952 241486 137964
rect 385678 137952 385684 137964
rect 241480 137924 385684 137952
rect 241480 137912 241486 137924
rect 385678 137912 385684 137924
rect 385736 137912 385742 137964
rect 35342 135124 35348 135176
rect 35400 135164 35406 135176
rect 38010 135164 38016 135176
rect 35400 135136 38016 135164
rect 35400 135124 35406 135136
rect 38010 135124 38016 135136
rect 38068 135124 38074 135176
rect 38286 128324 38292 128376
rect 38344 128364 38350 128376
rect 40494 128364 40500 128376
rect 38344 128336 40500 128364
rect 38344 128324 38350 128336
rect 40494 128324 40500 128336
rect 40552 128324 40558 128376
rect 241422 128256 241428 128308
rect 241480 128296 241486 128308
rect 294598 128296 294604 128308
rect 241480 128268 294604 128296
rect 241480 128256 241486 128268
rect 294598 128256 294604 128268
rect 294656 128256 294662 128308
rect 341518 126896 341524 126948
rect 341576 126936 341582 126948
rect 580166 126936 580172 126948
rect 341576 126908 580172 126936
rect 341576 126896 341582 126908
rect 580166 126896 580172 126908
rect 580224 126896 580230 126948
rect 35710 124108 35716 124160
rect 35768 124148 35774 124160
rect 38010 124148 38016 124160
rect 35768 124120 38016 124148
rect 35768 124108 35774 124120
rect 38010 124108 38016 124120
rect 38068 124108 38074 124160
rect 279418 113092 279424 113144
rect 279476 113132 279482 113144
rect 579614 113132 579620 113144
rect 279476 113104 579620 113132
rect 279476 113092 279482 113104
rect 579614 113092 579620 113104
rect 579672 113092 579678 113144
rect 240870 113024 240876 113076
rect 240928 113064 240934 113076
rect 291838 113064 291844 113076
rect 240928 113036 291844 113064
rect 240928 113024 240934 113036
rect 291838 113024 291844 113036
rect 291896 113024 291902 113076
rect 3142 111732 3148 111784
rect 3200 111772 3206 111784
rect 19978 111772 19984 111784
rect 3200 111744 19984 111772
rect 3200 111732 3206 111744
rect 19978 111732 19984 111744
rect 20036 111732 20042 111784
rect 35434 107584 35440 107636
rect 35492 107624 35498 107636
rect 38010 107624 38016 107636
rect 35492 107596 38016 107624
rect 35492 107584 35498 107596
rect 38010 107584 38016 107596
rect 38068 107584 38074 107636
rect 241422 107584 241428 107636
rect 241480 107624 241486 107636
rect 367738 107624 367744 107636
rect 241480 107596 367744 107624
rect 241480 107584 241486 107596
rect 367738 107584 367744 107596
rect 367796 107584 367802 107636
rect 241238 103436 241244 103488
rect 241296 103476 241302 103488
rect 337470 103476 337476 103488
rect 241296 103448 337476 103476
rect 241296 103436 241302 103448
rect 337470 103436 337476 103448
rect 337528 103436 337534 103488
rect 283558 100648 283564 100700
rect 283616 100688 283622 100700
rect 580166 100688 580172 100700
rect 283616 100660 580172 100688
rect 283616 100648 283622 100660
rect 580166 100648 580172 100660
rect 580224 100648 580230 100700
rect 241422 93780 241428 93832
rect 241480 93820 241486 93832
rect 373258 93820 373264 93832
rect 241480 93792 373264 93820
rect 241480 93780 241486 93792
rect 373258 93780 373264 93792
rect 373316 93780 373322 93832
rect 241422 88272 241428 88324
rect 241480 88312 241486 88324
rect 361574 88312 361580 88324
rect 241480 88284 361580 88312
rect 241480 88272 241486 88284
rect 361574 88272 361580 88284
rect 361632 88272 361638 88324
rect 268378 86912 268384 86964
rect 268436 86952 268442 86964
rect 579614 86952 579620 86964
rect 268436 86924 579620 86952
rect 268436 86912 268442 86924
rect 579614 86912 579620 86924
rect 579672 86912 579678 86964
rect 3142 85484 3148 85536
rect 3200 85524 3206 85536
rect 25498 85524 25504 85536
rect 3200 85496 25504 85524
rect 3200 85484 3206 85496
rect 25498 85484 25504 85496
rect 25556 85484 25562 85536
rect 241238 78616 241244 78668
rect 241296 78656 241302 78668
rect 360194 78656 360200 78668
rect 241296 78628 360200 78656
rect 241296 78616 241302 78628
rect 360194 78616 360200 78628
rect 360252 78616 360258 78668
rect 35526 75828 35532 75880
rect 35584 75868 35590 75880
rect 38010 75868 38016 75880
rect 35584 75840 38016 75868
rect 35584 75828 35590 75840
rect 38010 75828 38016 75840
rect 38068 75828 38074 75880
rect 276658 73108 276664 73160
rect 276716 73148 276722 73160
rect 580166 73148 580172 73160
rect 276716 73120 580172 73148
rect 276716 73108 276722 73120
rect 580166 73108 580172 73120
rect 580224 73108 580230 73160
rect 3142 71612 3148 71664
rect 3200 71652 3206 71664
rect 6178 71652 6184 71664
rect 3200 71624 6184 71652
rect 3200 71612 3206 71624
rect 6178 71612 6184 71624
rect 6236 71612 6242 71664
rect 241422 67532 241428 67584
rect 241480 67572 241486 67584
rect 351178 67572 351184 67584
rect 241480 67544 351184 67572
rect 241480 67532 241486 67544
rect 351178 67532 351184 67544
rect 351236 67532 351242 67584
rect 241238 63452 241244 63504
rect 241296 63492 241302 63504
rect 358814 63492 358820 63504
rect 241296 63464 358820 63492
rect 241296 63452 241302 63464
rect 358814 63452 358820 63464
rect 358872 63452 358878 63504
rect 3050 59304 3056 59356
rect 3108 59344 3114 59356
rect 13078 59344 13084 59356
rect 3108 59316 13084 59344
rect 3108 59304 3114 59316
rect 13078 59304 13084 59316
rect 13136 59304 13142 59356
rect 241422 52368 241428 52420
rect 241480 52408 241486 52420
rect 362954 52408 362960 52420
rect 241480 52380 362960 52408
rect 241480 52368 241486 52380
rect 362954 52368 362960 52380
rect 363012 52368 363018 52420
rect 266998 46860 267004 46912
rect 267056 46900 267062 46912
rect 580166 46900 580172 46912
rect 267056 46872 580172 46900
rect 267056 46860 267062 46872
rect 580166 46860 580172 46872
rect 580224 46860 580230 46912
rect 3418 45500 3424 45552
rect 3476 45540 3482 45552
rect 28258 45540 28264 45552
rect 3476 45512 28264 45540
rect 3476 45500 3482 45512
rect 28258 45500 28264 45512
rect 28316 45500 28322 45552
rect 35802 42712 35808 42764
rect 35860 42752 35866 42764
rect 38010 42752 38016 42764
rect 35860 42724 38016 42752
rect 35860 42712 35866 42724
rect 38010 42712 38016 42724
rect 38068 42712 38074 42764
rect 58268 40072 191604 40100
rect 58268 39908 58296 40072
rect 191576 39908 191604 40072
rect 58250 39856 58256 39908
rect 58308 39856 58314 39908
rect 191558 39856 191564 39908
rect 191616 39856 191622 39908
rect 234890 39856 234896 39908
rect 234948 39896 234954 39908
rect 238846 39896 238852 39908
rect 234948 39868 238852 39896
rect 234948 39856 234954 39868
rect 238846 39856 238852 39868
rect 238904 39856 238910 39908
rect 233510 39380 233516 39432
rect 233568 39420 233574 39432
rect 241514 39420 241520 39432
rect 233568 39392 241520 39420
rect 233568 39380 233574 39392
rect 241514 39380 241520 39392
rect 241572 39380 241578 39432
rect 38470 39312 38476 39364
rect 38528 39352 38534 39364
rect 106458 39352 106464 39364
rect 38528 39324 106464 39352
rect 38528 39312 38534 39324
rect 106458 39312 106464 39324
rect 106516 39312 106522 39364
rect 202046 39312 202052 39364
rect 202104 39352 202110 39364
rect 255958 39352 255964 39364
rect 202104 39324 255964 39352
rect 202104 39312 202110 39324
rect 255958 39312 255964 39324
rect 256016 39312 256022 39364
rect 196802 39244 196808 39296
rect 196860 39284 196866 39296
rect 287698 39284 287704 39296
rect 196860 39256 287704 39284
rect 196860 39244 196866 39256
rect 287698 39244 287704 39256
rect 287756 39244 287762 39296
rect 199470 39176 199476 39228
rect 199528 39216 199534 39228
rect 352558 39216 352564 39228
rect 199528 39188 352564 39216
rect 199528 39176 199534 39188
rect 352558 39176 352564 39188
rect 352616 39176 352622 39228
rect 232222 39108 232228 39160
rect 232280 39148 232286 39160
rect 411898 39148 411904 39160
rect 232280 39120 411904 39148
rect 232280 39108 232286 39120
rect 411898 39108 411904 39120
rect 411956 39108 411962 39160
rect 223022 39040 223028 39092
rect 223080 39080 223086 39092
rect 406378 39080 406384 39092
rect 223080 39052 406384 39080
rect 223080 39040 223086 39052
rect 406378 39040 406384 39052
rect 406436 39040 406442 39092
rect 224402 38972 224408 39024
rect 224460 39012 224466 39024
rect 409138 39012 409144 39024
rect 224460 38984 409144 39012
rect 224460 38972 224466 38984
rect 409138 38972 409144 38984
rect 409196 38972 409202 39024
rect 211246 38904 211252 38956
rect 211304 38944 211310 38956
rect 399478 38944 399484 38956
rect 211304 38916 399484 38944
rect 211304 38904 211310 38916
rect 399478 38904 399484 38916
rect 399536 38904 399542 38956
rect 212534 38836 212540 38888
rect 212592 38876 212598 38888
rect 402238 38876 402244 38888
rect 212592 38848 402244 38876
rect 212592 38836 212598 38848
rect 402238 38836 402244 38848
rect 402296 38836 402302 38888
rect 206002 38768 206008 38820
rect 206060 38808 206066 38820
rect 395338 38808 395344 38820
rect 206060 38780 395344 38808
rect 206060 38768 206066 38780
rect 395338 38768 395344 38780
rect 395396 38768 395402 38820
rect 221734 38700 221740 38752
rect 221792 38740 221798 38752
rect 420914 38740 420920 38752
rect 221792 38712 420920 38740
rect 221792 38700 221798 38712
rect 420914 38700 420920 38712
rect 420972 38700 420978 38752
rect 228266 38632 228272 38684
rect 228324 38672 228330 38684
rect 434714 38672 434720 38684
rect 228324 38644 434720 38672
rect 228324 38632 228330 38644
rect 434714 38632 434720 38644
rect 434772 38632 434778 38684
rect 39298 38564 39304 38616
rect 39356 38604 39362 38616
rect 40678 38604 40684 38616
rect 39356 38576 40684 38604
rect 39356 38564 39362 38576
rect 40678 38564 40684 38576
rect 40736 38604 40742 38616
rect 183646 38604 183652 38616
rect 40736 38576 183652 38604
rect 40736 38564 40742 38576
rect 183646 38564 183652 38576
rect 183704 38564 183710 38616
rect 217778 38564 217784 38616
rect 217836 38604 217842 38616
rect 237926 38604 237932 38616
rect 217836 38576 237932 38604
rect 217836 38564 217842 38576
rect 237926 38564 237932 38576
rect 237984 38564 237990 38616
rect 40310 38496 40316 38548
rect 40368 38536 40374 38548
rect 186314 38536 186320 38548
rect 40368 38508 186320 38536
rect 40368 38496 40374 38508
rect 186314 38496 186320 38508
rect 186372 38496 186378 38548
rect 220446 38496 220452 38548
rect 220504 38536 220510 38548
rect 238110 38536 238116 38548
rect 220504 38508 238116 38536
rect 220504 38496 220510 38508
rect 238110 38496 238116 38508
rect 238168 38496 238174 38548
rect 51718 38428 51724 38480
rect 51776 38468 51782 38480
rect 61654 38468 61660 38480
rect 51776 38440 61660 38468
rect 51776 38428 51782 38440
rect 61654 38428 61660 38440
rect 61712 38428 61718 38480
rect 106458 38428 106464 38480
rect 106516 38468 106522 38480
rect 195514 38468 195520 38480
rect 106516 38440 195520 38468
rect 106516 38428 106522 38440
rect 195514 38428 195520 38440
rect 195572 38428 195578 38480
rect 229646 38428 229652 38480
rect 229704 38468 229710 38480
rect 392578 38468 392584 38480
rect 229704 38440 392584 38468
rect 229704 38428 229710 38440
rect 392578 38428 392584 38440
rect 392636 38428 392642 38480
rect 53098 38360 53104 38412
rect 53156 38400 53162 38412
rect 87874 38400 87880 38412
rect 53156 38372 87880 38400
rect 53156 38360 53162 38372
rect 87874 38360 87880 38372
rect 87932 38360 87938 38412
rect 226978 38360 226984 38412
rect 227036 38400 227042 38412
rect 238018 38400 238024 38412
rect 227036 38372 238024 38400
rect 227036 38360 227042 38372
rect 238018 38360 238024 38372
rect 238076 38360 238082 38412
rect 10962 38292 10968 38344
rect 11020 38332 11026 38344
rect 51166 38332 51172 38344
rect 11020 38304 51172 38332
rect 11020 38292 11026 38304
rect 51166 38292 51172 38304
rect 51224 38292 51230 38344
rect 54478 38292 54484 38344
rect 54536 38332 54542 38344
rect 91830 38332 91836 38344
rect 54536 38304 91836 38332
rect 54536 38292 54542 38304
rect 91830 38292 91836 38304
rect 91888 38292 91894 38344
rect 190270 38292 190276 38344
rect 190328 38332 190334 38344
rect 258718 38332 258724 38344
rect 190328 38304 258724 38332
rect 190328 38292 190334 38304
rect 258718 38292 258724 38304
rect 258776 38292 258782 38344
rect 15102 38224 15108 38276
rect 15160 38264 15166 38276
rect 56410 38264 56416 38276
rect 15160 38236 56416 38264
rect 15160 38224 15166 38236
rect 56410 38224 56416 38236
rect 56468 38224 56474 38276
rect 60366 38224 60372 38276
rect 60424 38264 60430 38276
rect 68186 38264 68192 38276
rect 60424 38236 68192 38264
rect 60424 38224 60430 38236
rect 68186 38224 68192 38236
rect 68244 38224 68250 38276
rect 194134 38224 194140 38276
rect 194192 38264 194198 38276
rect 261478 38264 261484 38276
rect 194192 38236 261484 38264
rect 194192 38224 194198 38236
rect 261478 38224 261484 38236
rect 261536 38224 261542 38276
rect 24762 38156 24768 38208
rect 24820 38196 24826 38208
rect 66898 38196 66904 38208
rect 24820 38168 66904 38196
rect 24820 38156 24826 38168
rect 66898 38156 66904 38168
rect 66956 38156 66962 38208
rect 198090 38156 198096 38208
rect 198148 38196 198154 38208
rect 262858 38196 262864 38208
rect 198148 38168 262864 38196
rect 198148 38156 198154 38168
rect 262858 38156 262864 38168
rect 262916 38156 262922 38208
rect 37182 38088 37188 38140
rect 37240 38128 37246 38140
rect 79962 38128 79968 38140
rect 37240 38100 79968 38128
rect 37240 38088 37246 38100
rect 79962 38088 79968 38100
rect 80020 38088 80026 38140
rect 225690 38088 225696 38140
rect 225748 38128 225754 38140
rect 290458 38128 290464 38140
rect 225748 38100 290464 38128
rect 225748 38088 225754 38100
rect 290458 38088 290464 38100
rect 290516 38088 290522 38140
rect 33042 38020 33048 38072
rect 33100 38060 33106 38072
rect 76098 38060 76104 38072
rect 33100 38032 76104 38060
rect 33100 38020 33106 38032
rect 76098 38020 76104 38032
rect 76156 38020 76162 38072
rect 208578 38020 208584 38072
rect 208636 38060 208642 38072
rect 250438 38060 250444 38072
rect 208636 38032 250444 38060
rect 208636 38020 208642 38032
rect 250438 38020 250444 38032
rect 250496 38020 250502 38072
rect 28902 37952 28908 38004
rect 28960 37992 28966 38004
rect 72142 37992 72148 38004
rect 28960 37964 72148 37992
rect 28960 37952 28966 37964
rect 72142 37952 72148 37964
rect 72200 37952 72206 38004
rect 81434 37952 81440 38004
rect 81492 37992 81498 38004
rect 82630 37992 82636 38004
rect 81492 37964 82636 37992
rect 81492 37952 81498 37964
rect 82630 37952 82636 37964
rect 82688 37952 82694 38004
rect 106366 37952 106372 38004
rect 106424 37992 106430 38004
rect 107562 37992 107568 38004
rect 106424 37964 107568 37992
rect 106424 37952 106430 37964
rect 107562 37952 107568 37964
rect 107620 37952 107626 38004
rect 135254 37952 135260 38004
rect 135312 37992 135318 38004
rect 136450 37992 136456 38004
rect 135312 37964 136456 37992
rect 135312 37952 135318 37964
rect 136450 37952 136456 37964
rect 136508 37952 136514 38004
rect 159358 37952 159364 38004
rect 159416 37992 159422 38004
rect 160094 37992 160100 38004
rect 159416 37964 160100 37992
rect 159416 37952 159422 37964
rect 160094 37952 160100 37964
rect 160152 37952 160158 38004
rect 160186 37952 160192 38004
rect 160244 37992 160250 38004
rect 161382 37992 161388 38004
rect 160244 37964 161388 37992
rect 160244 37952 160250 37964
rect 161382 37952 161388 37964
rect 161440 37952 161446 38004
rect 161474 37952 161480 38004
rect 161532 37992 161538 38004
rect 162670 37992 162676 38004
rect 161532 37964 162676 37992
rect 161532 37952 161538 37964
rect 162670 37952 162676 37964
rect 162728 37952 162734 38004
rect 179782 37952 179788 38004
rect 179840 37992 179846 38004
rect 180702 37992 180708 38004
rect 179840 37964 180708 37992
rect 179840 37952 179846 37964
rect 180702 37952 180708 37964
rect 180760 37952 180766 38004
rect 182358 37952 182364 38004
rect 182416 37992 182422 38004
rect 183462 37992 183468 38004
rect 182416 37964 183468 37992
rect 182416 37952 182422 37964
rect 183462 37952 183468 37964
rect 183520 37952 183526 38004
rect 213822 37952 213828 38004
rect 213880 37992 213886 38004
rect 380158 37992 380164 38004
rect 213880 37964 380164 37992
rect 213880 37952 213886 37964
rect 380158 37952 380164 37964
rect 380216 37952 380222 38004
rect 39942 37884 39948 37936
rect 40000 37924 40006 37936
rect 83918 37924 83924 37936
rect 40000 37896 83924 37924
rect 40000 37884 40006 37896
rect 83918 37884 83924 37896
rect 83976 37884 83982 37936
rect 162118 37884 162124 37936
rect 162176 37924 162182 37936
rect 163958 37924 163964 37936
rect 162176 37896 163964 37924
rect 162176 37884 162182 37896
rect 163958 37884 163964 37896
rect 164016 37884 164022 37936
rect 219158 37884 219164 37936
rect 219216 37924 219222 37936
rect 384298 37924 384304 37936
rect 219216 37896 384304 37924
rect 219216 37884 219222 37896
rect 384298 37884 384304 37896
rect 384356 37884 384362 37936
rect 55858 37816 55864 37868
rect 55916 37856 55922 37868
rect 57698 37856 57704 37868
rect 55916 37828 57704 37856
rect 55916 37816 55922 37828
rect 57698 37816 57704 37828
rect 57756 37816 57762 37868
rect 100018 37816 100024 37868
rect 100076 37856 100082 37868
rect 101030 37856 101036 37868
rect 100076 37828 101036 37856
rect 100076 37816 100082 37828
rect 101030 37816 101036 37828
rect 101088 37816 101094 37868
rect 181070 37816 181076 37868
rect 181128 37856 181134 37868
rect 182082 37856 182088 37868
rect 181128 37828 182088 37856
rect 181128 37816 181134 37828
rect 182082 37816 182088 37828
rect 182140 37816 182146 37868
rect 185026 37748 185032 37800
rect 185084 37788 185090 37800
rect 254578 37788 254584 37800
rect 185084 37760 254584 37788
rect 185084 37748 185090 37760
rect 254578 37748 254584 37760
rect 254636 37748 254642 37800
rect 57238 37680 57244 37732
rect 57296 37720 57302 37732
rect 62942 37720 62948 37732
rect 57296 37692 62948 37720
rect 57296 37680 57302 37692
rect 62942 37680 62948 37692
rect 63000 37680 63006 37732
rect 95878 37680 95884 37732
rect 95936 37720 95942 37732
rect 99650 37720 99656 37732
rect 95936 37692 99656 37720
rect 95936 37680 95942 37692
rect 99650 37680 99656 37692
rect 99708 37680 99714 37732
rect 209958 37680 209964 37732
rect 210016 37720 210022 37732
rect 238202 37720 238208 37732
rect 210016 37692 238208 37720
rect 210016 37680 210022 37692
rect 238202 37680 238208 37692
rect 238260 37680 238266 37732
rect 230934 37612 230940 37664
rect 230992 37652 230998 37664
rect 239030 37652 239036 37664
rect 230992 37624 239036 37652
rect 230992 37612 230998 37624
rect 239030 37612 239036 37624
rect 239088 37612 239094 37664
rect 236178 37544 236184 37596
rect 236236 37584 236242 37596
rect 241606 37584 241612 37596
rect 236236 37556 241612 37584
rect 236236 37544 236242 37556
rect 241606 37544 241612 37556
rect 241664 37544 241670 37596
rect 91738 37272 91744 37324
rect 91796 37312 91802 37324
rect 94406 37312 94412 37324
rect 91796 37284 94412 37312
rect 91796 37272 91802 37284
rect 94406 37272 94412 37284
rect 94464 37272 94470 37324
rect 151078 37272 151084 37324
rect 151136 37312 151142 37324
rect 152182 37312 152188 37324
rect 151136 37284 152188 37312
rect 151136 37272 151142 37284
rect 152182 37272 152188 37284
rect 152240 37272 152246 37324
rect 72418 37204 72424 37256
rect 72476 37244 72482 37256
rect 110230 37244 110236 37256
rect 72476 37216 110236 37244
rect 72476 37204 72482 37216
rect 110230 37204 110236 37216
rect 110288 37204 110294 37256
rect 25498 37136 25504 37188
rect 25556 37176 25562 37188
rect 49786 37176 49792 37188
rect 25556 37148 49792 37176
rect 25556 37136 25562 37148
rect 49786 37136 49792 37148
rect 49844 37136 49850 37188
rect 75178 37136 75184 37188
rect 75236 37176 75242 37188
rect 114094 37176 114100 37188
rect 75236 37148 114100 37176
rect 75236 37136 75242 37148
rect 114094 37136 114100 37148
rect 114152 37136 114158 37188
rect 15838 37068 15844 37120
rect 15896 37108 15902 37120
rect 43254 37108 43260 37120
rect 15896 37080 43260 37108
rect 15896 37068 15902 37080
rect 43254 37068 43260 37080
rect 43312 37068 43318 37120
rect 90358 37068 90364 37120
rect 90416 37108 90422 37120
rect 135162 37108 135168 37120
rect 90416 37080 135168 37108
rect 90416 37068 90422 37080
rect 135162 37068 135168 37080
rect 135220 37068 135226 37120
rect 6178 37000 6184 37052
rect 6236 37040 6242 37052
rect 38562 37040 38568 37052
rect 6236 37012 38568 37040
rect 6236 37000 6242 37012
rect 38562 37000 38568 37012
rect 38620 37040 38626 37052
rect 41966 37040 41972 37052
rect 38620 37012 41972 37040
rect 38620 37000 38626 37012
rect 41966 37000 41972 37012
rect 42024 37000 42030 37052
rect 43438 37000 43444 37052
rect 43496 37040 43502 37052
rect 69474 37040 69480 37052
rect 43496 37012 69480 37040
rect 43496 37000 43502 37012
rect 69474 37000 69480 37012
rect 69532 37000 69538 37052
rect 87598 37000 87604 37052
rect 87656 37040 87662 37052
rect 131206 37040 131212 37052
rect 87656 37012 131212 37040
rect 87656 37000 87662 37012
rect 131206 37000 131212 37012
rect 131264 37000 131270 37052
rect 17218 36932 17224 36984
rect 17276 36972 17282 36984
rect 53742 36972 53748 36984
rect 17276 36944 53748 36972
rect 17276 36932 17282 36944
rect 53742 36932 53748 36944
rect 53800 36932 53806 36984
rect 70302 36932 70308 36984
rect 70360 36972 70366 36984
rect 116762 36972 116768 36984
rect 70360 36944 116768 36972
rect 70360 36932 70366 36944
rect 116762 36932 116768 36944
rect 116820 36932 116826 36984
rect 19978 36864 19984 36916
rect 20036 36904 20042 36916
rect 58986 36904 58992 36916
rect 20036 36876 58992 36904
rect 20036 36864 20042 36876
rect 58986 36864 58992 36876
rect 59044 36864 59050 36916
rect 66162 36864 66168 36916
rect 66220 36904 66226 36916
rect 112806 36904 112812 36916
rect 66220 36876 112812 36904
rect 66220 36864 66226 36876
rect 112806 36864 112812 36876
rect 112864 36864 112870 36916
rect 131758 36864 131764 36916
rect 131816 36904 131822 36916
rect 145650 36904 145656 36916
rect 131816 36876 145656 36904
rect 131816 36864 131822 36876
rect 145650 36864 145656 36876
rect 145708 36864 145714 36916
rect 4062 36796 4068 36848
rect 4120 36836 4126 36848
rect 44542 36836 44548 36848
rect 4120 36808 44548 36836
rect 4120 36796 4126 36808
rect 44542 36796 44548 36808
rect 44600 36796 44606 36848
rect 48958 36796 48964 36848
rect 49016 36836 49022 36848
rect 81342 36836 81348 36848
rect 49016 36808 81348 36836
rect 49016 36796 49022 36808
rect 81342 36796 81348 36808
rect 81400 36796 81406 36848
rect 86218 36796 86224 36848
rect 86276 36836 86282 36848
rect 133782 36836 133788 36848
rect 86276 36808 133788 36836
rect 86276 36796 86282 36808
rect 133782 36796 133788 36808
rect 133840 36796 133846 36848
rect 142798 36796 142804 36848
rect 142856 36836 142862 36848
rect 173158 36836 173164 36848
rect 142856 36808 173164 36836
rect 142856 36796 142862 36808
rect 173158 36796 173164 36808
rect 173216 36796 173222 36848
rect 13722 36728 13728 36780
rect 13780 36768 13786 36780
rect 55030 36768 55036 36780
rect 13780 36740 55036 36768
rect 13780 36728 13786 36740
rect 55030 36728 55036 36740
rect 55088 36728 55094 36780
rect 66898 36728 66904 36780
rect 66956 36768 66962 36780
rect 98362 36768 98368 36780
rect 66956 36740 98368 36768
rect 66956 36728 66962 36740
rect 98362 36728 98368 36740
rect 98420 36728 98426 36780
rect 101398 36728 101404 36780
rect 101456 36768 101462 36780
rect 150894 36768 150900 36780
rect 101456 36740 150900 36768
rect 101456 36728 101462 36740
rect 150894 36728 150900 36740
rect 150952 36728 150958 36780
rect 31662 36660 31668 36712
rect 31720 36700 31726 36712
rect 74718 36700 74724 36712
rect 31720 36672 74724 36700
rect 31720 36660 31726 36672
rect 74718 36660 74724 36672
rect 74776 36660 74782 36712
rect 83458 36660 83464 36712
rect 83516 36700 83522 36712
rect 90542 36700 90548 36712
rect 83516 36672 90548 36700
rect 83516 36660 83522 36672
rect 90542 36660 90548 36672
rect 90600 36660 90606 36712
rect 108298 36660 108304 36712
rect 108356 36700 108362 36712
rect 158714 36700 158720 36712
rect 108356 36672 158720 36700
rect 108356 36660 108362 36672
rect 158714 36660 158720 36672
rect 158772 36660 158778 36712
rect 8202 36592 8208 36644
rect 8260 36632 8266 36644
rect 48498 36632 48504 36644
rect 8260 36604 48504 36632
rect 8260 36592 8266 36604
rect 48498 36592 48504 36604
rect 48556 36592 48562 36644
rect 62022 36592 62028 36644
rect 62080 36632 62086 36644
rect 108850 36632 108856 36644
rect 62080 36604 108856 36632
rect 62080 36592 62086 36604
rect 108850 36592 108856 36604
rect 108908 36592 108914 36644
rect 114462 36592 114468 36644
rect 114520 36632 114526 36644
rect 166626 36632 166632 36644
rect 114520 36604 166632 36632
rect 114520 36592 114526 36604
rect 166626 36592 166632 36604
rect 166684 36592 166690 36644
rect 2038 36524 2044 36576
rect 2096 36564 2102 36576
rect 40678 36564 40684 36576
rect 2096 36536 40684 36564
rect 2096 36524 2102 36536
rect 40678 36524 40684 36536
rect 40736 36524 40742 36576
rect 42702 36524 42708 36576
rect 42760 36564 42766 36576
rect 86586 36564 86592 36576
rect 42760 36536 86592 36564
rect 42760 36524 42766 36536
rect 86586 36524 86592 36536
rect 86644 36524 86650 36576
rect 104802 36524 104808 36576
rect 104860 36564 104866 36576
rect 156138 36564 156144 36576
rect 104860 36536 156144 36564
rect 104860 36524 104866 36536
rect 156138 36524 156144 36536
rect 156196 36524 156202 36576
rect 71038 36456 71044 36508
rect 71096 36496 71102 36508
rect 106274 36496 106280 36508
rect 71096 36468 106280 36496
rect 71096 36456 71102 36468
rect 106274 36456 106280 36468
rect 106332 36456 106338 36508
rect 68278 36388 68284 36440
rect 68336 36428 68342 36440
rect 102318 36428 102324 36440
rect 68336 36400 102324 36428
rect 68336 36388 68342 36400
rect 102318 36388 102324 36400
rect 102376 36388 102382 36440
rect 50982 35164 50988 35216
rect 51040 35204 51046 35216
rect 95786 35204 95792 35216
rect 51040 35176 95792 35204
rect 51040 35164 51046 35176
rect 95786 35164 95792 35176
rect 95844 35164 95850 35216
rect 2866 33056 2872 33108
rect 2924 33096 2930 33108
rect 21358 33096 21364 33108
rect 2924 33068 21364 33096
rect 2924 33056 2930 33068
rect 21358 33056 21364 33068
rect 21416 33056 21422 33108
rect 273898 33056 273904 33108
rect 273956 33096 273962 33108
rect 580166 33096 580172 33108
rect 273956 33068 580172 33096
rect 273956 33056 273962 33068
rect 580166 33056 580172 33068
rect 580224 33056 580230 33108
rect 21450 32376 21456 32428
rect 21508 32416 21514 32428
rect 59354 32416 59360 32428
rect 21508 32388 59360 32416
rect 21508 32376 21514 32388
rect 59354 32376 59360 32388
rect 59412 32376 59418 32428
rect 3418 20612 3424 20664
rect 3476 20652 3482 20664
rect 14458 20652 14464 20664
rect 3476 20624 14464 20652
rect 3476 20612 3482 20624
rect 14458 20612 14464 20624
rect 14516 20612 14522 20664
rect 111610 11772 111616 11824
rect 111668 11812 111674 11824
rect 162118 11812 162124 11824
rect 111668 11784 162124 11812
rect 111668 11772 111674 11784
rect 162118 11772 162124 11784
rect 162176 11772 162182 11824
rect 33870 11704 33876 11756
rect 33928 11744 33934 11756
rect 64874 11744 64880 11756
rect 33928 11716 64880 11744
rect 33928 11704 33934 11716
rect 64874 11704 64880 11716
rect 64932 11704 64938 11756
rect 115842 11704 115848 11756
rect 115900 11744 115906 11756
rect 166994 11744 167000 11756
rect 115900 11716 167000 11744
rect 115900 11704 115906 11716
rect 166994 11704 167000 11716
rect 167052 11704 167058 11756
rect 105538 10276 105544 10328
rect 105596 10316 105602 10328
rect 142154 10316 142160 10328
rect 105596 10288 142160 10316
rect 105596 10276 105602 10288
rect 142154 10276 142160 10288
rect 142212 10276 142218 10328
rect 61930 7556 61936 7608
rect 61988 7596 61994 7608
rect 104894 7596 104900 7608
rect 61988 7568 104900 7596
rect 61988 7556 61994 7568
rect 104894 7556 104900 7568
rect 104952 7556 104958 7608
rect 3418 6808 3424 6860
rect 3476 6848 3482 6860
rect 33778 6848 33784 6860
rect 3476 6820 33784 6848
rect 3476 6808 3482 6820
rect 33778 6808 33784 6820
rect 33836 6808 33842 6860
rect 265618 6808 265624 6860
rect 265676 6848 265682 6860
rect 580166 6848 580172 6860
rect 265676 6820 580172 6848
rect 265676 6808 265682 6820
rect 580166 6808 580172 6820
rect 580224 6808 580230 6860
rect 92566 6604 92572 6656
rect 92624 6644 92630 6656
rect 125594 6644 125600 6656
rect 92624 6616 125600 6644
rect 92624 6604 92630 6616
rect 125594 6604 125600 6616
rect 125652 6604 125658 6656
rect 87506 6536 87512 6588
rect 87564 6576 87570 6588
rect 117314 6576 117320 6588
rect 87564 6548 117320 6576
rect 87564 6536 87570 6548
rect 117314 6536 117320 6548
rect 117372 6536 117378 6588
rect 117958 6536 117964 6588
rect 118016 6576 118022 6588
rect 153194 6576 153200 6588
rect 118016 6548 153200 6576
rect 118016 6536 118022 6548
rect 153194 6536 153200 6548
rect 153252 6536 153258 6588
rect 99374 6468 99380 6520
rect 99432 6508 99438 6520
rect 140774 6508 140780 6520
rect 99432 6480 140780 6508
rect 99432 6468 99438 6480
rect 140774 6468 140780 6480
rect 140832 6468 140838 6520
rect 38378 6400 38384 6452
rect 38436 6440 38442 6452
rect 81434 6440 81440 6452
rect 38436 6412 81440 6440
rect 38436 6400 38442 6412
rect 81434 6400 81440 6412
rect 81492 6400 81498 6452
rect 88426 6400 88432 6452
rect 88484 6440 88490 6452
rect 136634 6440 136640 6452
rect 88484 6412 136640 6440
rect 88484 6400 88490 6412
rect 136634 6400 136640 6412
rect 136692 6400 136698 6452
rect 47854 6332 47860 6384
rect 47912 6372 47918 6384
rect 92474 6372 92480 6384
rect 47912 6344 92480 6372
rect 47912 6332 47918 6344
rect 92474 6332 92480 6344
rect 92532 6332 92538 6384
rect 101030 6332 101036 6384
rect 101088 6372 101094 6384
rect 151078 6372 151084 6384
rect 101088 6344 151084 6372
rect 101088 6332 101094 6344
rect 151078 6332 151084 6344
rect 151136 6332 151142 6384
rect 51350 6264 51356 6316
rect 51408 6304 51414 6316
rect 96614 6304 96620 6316
rect 51408 6276 96620 6304
rect 51408 6264 51414 6276
rect 96614 6264 96620 6276
rect 96672 6264 96678 6316
rect 108114 6264 108120 6316
rect 108172 6304 108178 6316
rect 159358 6304 159364 6316
rect 108172 6276 159364 6304
rect 108172 6264 108178 6276
rect 159358 6264 159364 6276
rect 159416 6264 159422 6316
rect 54938 6196 54944 6248
rect 54996 6236 55002 6248
rect 100018 6236 100024 6248
rect 54996 6208 100024 6236
rect 54996 6196 55002 6208
rect 100018 6196 100024 6208
rect 100076 6196 100082 6248
rect 118786 6196 118792 6248
rect 118844 6236 118850 6248
rect 171134 6236 171140 6248
rect 118844 6208 171140 6236
rect 118844 6196 118850 6208
rect 171134 6196 171140 6208
rect 171192 6196 171198 6248
rect 73798 6128 73804 6180
rect 73856 6168 73862 6180
rect 121454 6168 121460 6180
rect 73856 6140 121460 6168
rect 73856 6128 73862 6140
rect 121454 6128 121460 6140
rect 121512 6128 121518 6180
rect 122282 6128 122288 6180
rect 122340 6168 122346 6180
rect 175274 6168 175280 6180
rect 122340 6140 175280 6168
rect 122340 6128 122346 6140
rect 175274 6128 175280 6140
rect 175332 6128 175338 6180
rect 83274 5448 83280 5500
rect 83332 5488 83338 5500
rect 132586 5488 132592 5500
rect 83332 5460 132592 5488
rect 83332 5448 83338 5460
rect 132586 5448 132592 5460
rect 132644 5448 132650 5500
rect 80882 5380 80888 5432
rect 80940 5420 80946 5432
rect 129734 5420 129740 5432
rect 80940 5392 129740 5420
rect 80940 5380 80946 5392
rect 129734 5380 129740 5392
rect 129792 5380 129798 5432
rect 79686 5312 79692 5364
rect 79744 5352 79750 5364
rect 128354 5352 128360 5364
rect 79744 5324 128360 5352
rect 79744 5312 79750 5324
rect 128354 5312 128360 5324
rect 128412 5312 128418 5364
rect 86862 5244 86868 5296
rect 86920 5284 86926 5296
rect 135254 5284 135260 5296
rect 86920 5256 135260 5284
rect 86920 5244 86926 5256
rect 135254 5244 135260 5256
rect 135312 5244 135318 5296
rect 51074 5176 51080 5228
rect 51132 5216 51138 5228
rect 88334 5216 88340 5228
rect 51132 5188 88340 5216
rect 51132 5176 51138 5188
rect 88334 5176 88340 5188
rect 88392 5176 88398 5228
rect 90358 5176 90364 5228
rect 90416 5216 90422 5228
rect 139394 5216 139400 5228
rect 90416 5188 139400 5216
rect 90416 5176 90422 5188
rect 139394 5176 139400 5188
rect 139452 5176 139458 5228
rect 49050 5108 49056 5160
rect 49108 5148 49114 5160
rect 91738 5148 91744 5160
rect 49108 5120 91744 5148
rect 49108 5108 49114 5120
rect 91738 5108 91744 5120
rect 91796 5108 91802 5160
rect 93946 5108 93952 5160
rect 94004 5148 94010 5160
rect 143534 5148 143540 5160
rect 94004 5120 143540 5148
rect 94004 5108 94010 5120
rect 143534 5108 143540 5120
rect 143592 5108 143598 5160
rect 40126 5040 40132 5092
rect 40184 5080 40190 5092
rect 77294 5080 77300 5092
rect 40184 5052 77300 5080
rect 40184 5040 40190 5052
rect 77294 5040 77300 5052
rect 77352 5040 77358 5092
rect 78582 5040 78588 5092
rect 78640 5080 78646 5092
rect 126974 5080 126980 5092
rect 78640 5052 126980 5080
rect 78640 5040 78646 5052
rect 126974 5040 126980 5052
rect 127032 5040 127038 5092
rect 128538 5040 128544 5092
rect 128596 5080 128602 5092
rect 178034 5080 178040 5092
rect 128596 5052 178040 5080
rect 128596 5040 128602 5052
rect 178034 5040 178040 5052
rect 178092 5040 178098 5092
rect 40678 4972 40684 5024
rect 40736 5012 40742 5024
rect 84194 5012 84200 5024
rect 40736 4984 84200 5012
rect 40736 4972 40742 4984
rect 84194 4972 84200 4984
rect 84252 4972 84258 5024
rect 98638 4972 98644 5024
rect 98696 5012 98702 5024
rect 149054 5012 149060 5024
rect 98696 4984 149060 5012
rect 98696 4972 98702 4984
rect 149054 4972 149060 4984
rect 149112 4972 149118 5024
rect 34790 4904 34796 4956
rect 34848 4944 34854 4956
rect 78766 4944 78772 4956
rect 34848 4916 78772 4944
rect 34848 4904 34854 4916
rect 78766 4904 78772 4916
rect 78824 4904 78830 4956
rect 97442 4904 97448 4956
rect 97500 4944 97506 4956
rect 147674 4944 147680 4956
rect 97500 4916 147680 4944
rect 97500 4904 97506 4916
rect 147674 4904 147680 4916
rect 147732 4904 147738 4956
rect 30098 4836 30104 4888
rect 30156 4876 30162 4888
rect 73154 4876 73160 4888
rect 30156 4848 73160 4876
rect 30156 4836 30162 4848
rect 73154 4836 73160 4848
rect 73212 4836 73218 4888
rect 105722 4836 105728 4888
rect 105780 4876 105786 4888
rect 157334 4876 157340 4888
rect 105780 4848 157340 4876
rect 105780 4836 105786 4848
rect 157334 4836 157340 4848
rect 157392 4836 157398 4888
rect 29822 4768 29828 4820
rect 29880 4808 29886 4820
rect 63402 4808 63408 4820
rect 29880 4780 63408 4808
rect 29880 4768 29886 4780
rect 63402 4768 63408 4780
rect 63460 4768 63466 4820
rect 63494 4768 63500 4820
rect 63552 4808 63558 4820
rect 70394 4808 70400 4820
rect 63552 4780 70400 4808
rect 63552 4768 63558 4780
rect 70394 4768 70400 4780
rect 70452 4768 70458 4820
rect 72602 4768 72608 4820
rect 72660 4808 72666 4820
rect 120074 4808 120080 4820
rect 72660 4780 120080 4808
rect 72660 4768 72666 4780
rect 120074 4768 120080 4780
rect 120132 4768 120138 4820
rect 123478 4768 123484 4820
rect 123536 4808 123542 4820
rect 176654 4808 176660 4820
rect 123536 4780 176660 4808
rect 123536 4768 123542 4780
rect 176654 4768 176660 4780
rect 176712 4768 176718 4820
rect 76190 4700 76196 4752
rect 76248 4740 76254 4752
rect 124214 4740 124220 4752
rect 76248 4712 124220 4740
rect 76248 4700 76254 4712
rect 124214 4700 124220 4712
rect 124272 4700 124278 4752
rect 74994 4632 75000 4684
rect 75052 4672 75058 4684
rect 122834 4672 122840 4684
rect 75052 4644 122840 4672
rect 75052 4632 75058 4644
rect 122834 4632 122840 4644
rect 122892 4632 122898 4684
rect 21818 4088 21824 4140
rect 21876 4128 21882 4140
rect 29822 4128 29828 4140
rect 21876 4100 29828 4128
rect 21876 4088 21882 4100
rect 29822 4088 29828 4100
rect 29880 4088 29886 4140
rect 43070 4088 43076 4140
rect 43128 4128 43134 4140
rect 53098 4128 53104 4140
rect 43128 4100 53104 4128
rect 43128 4088 43134 4100
rect 53098 4088 53104 4100
rect 53156 4088 53162 4140
rect 63218 4088 63224 4140
rect 63276 4128 63282 4140
rect 72418 4128 72424 4140
rect 63276 4100 72424 4128
rect 63276 4088 63282 4100
rect 72418 4088 72424 4100
rect 72476 4088 72482 4140
rect 91554 4088 91560 4140
rect 91612 4128 91618 4140
rect 99374 4128 99380 4140
rect 91612 4100 99380 4128
rect 91612 4088 91618 4100
rect 99374 4088 99380 4100
rect 99432 4088 99438 4140
rect 102226 4088 102232 4140
rect 102284 4128 102290 4140
rect 117958 4128 117964 4140
rect 102284 4100 117964 4128
rect 102284 4088 102290 4100
rect 117958 4088 117964 4100
rect 118016 4088 118022 4140
rect 119890 4088 119896 4140
rect 119948 4128 119954 4140
rect 142798 4128 142804 4140
rect 119948 4100 142804 4128
rect 119948 4088 119954 4100
rect 142798 4088 142804 4100
rect 142856 4088 142862 4140
rect 23014 4020 23020 4072
rect 23072 4060 23078 4072
rect 33870 4060 33876 4072
rect 23072 4032 33876 4060
rect 23072 4020 23078 4032
rect 33870 4020 33876 4032
rect 33928 4020 33934 4072
rect 37090 4020 37096 4072
rect 37148 4060 37154 4072
rect 48958 4060 48964 4072
rect 37148 4032 48964 4060
rect 37148 4020 37154 4032
rect 48958 4020 48964 4032
rect 49016 4020 49022 4072
rect 59630 4020 59636 4072
rect 59688 4060 59694 4072
rect 71038 4060 71044 4072
rect 59688 4032 71044 4060
rect 59688 4020 59694 4032
rect 71038 4020 71044 4032
rect 71096 4020 71102 4072
rect 77386 4020 77392 4072
rect 77444 4060 77450 4072
rect 92566 4060 92572 4072
rect 77444 4032 92572 4060
rect 77444 4020 77450 4032
rect 92566 4020 92572 4032
rect 92624 4020 92630 4072
rect 95142 4020 95148 4072
rect 95200 4060 95206 4072
rect 131758 4060 131764 4072
rect 95200 4032 131764 4060
rect 95200 4020 95206 4032
rect 131758 4020 131764 4032
rect 131816 4020 131822 4072
rect 19426 3952 19432 4004
rect 19484 3992 19490 4004
rect 51718 3992 51724 4004
rect 19484 3964 51724 3992
rect 19484 3952 19490 3964
rect 51718 3952 51724 3964
rect 51776 3952 51782 4004
rect 56042 3952 56048 4004
rect 56100 3992 56106 4004
rect 68278 3992 68284 4004
rect 56100 3964 68284 3992
rect 56100 3952 56106 3964
rect 68278 3952 68284 3964
rect 68336 3952 68342 4004
rect 82078 3952 82084 4004
rect 82136 3992 82142 4004
rect 87598 3992 87604 4004
rect 82136 3964 87604 3992
rect 82136 3952 82142 3964
rect 87598 3952 87604 3964
rect 87656 3952 87662 4004
rect 89162 3952 89168 4004
rect 89220 3992 89226 4004
rect 138014 3992 138020 4004
rect 89220 3964 138020 3992
rect 89220 3952 89226 3964
rect 138014 3952 138020 3964
rect 138072 3952 138078 4004
rect 27706 3884 27712 3936
rect 27764 3924 27770 3936
rect 63494 3924 63500 3936
rect 27764 3896 63500 3924
rect 27764 3884 27770 3896
rect 63494 3884 63500 3896
rect 63552 3884 63558 3936
rect 70210 3884 70216 3936
rect 70268 3924 70274 3936
rect 87506 3924 87512 3936
rect 70268 3896 87512 3924
rect 70268 3884 70274 3896
rect 87506 3884 87512 3896
rect 87564 3884 87570 3936
rect 92750 3884 92756 3936
rect 92808 3924 92814 3936
rect 105538 3924 105544 3936
rect 92808 3896 105544 3924
rect 92808 3884 92814 3896
rect 105538 3884 105544 3896
rect 105596 3884 105602 3936
rect 110506 3884 110512 3936
rect 110564 3924 110570 3936
rect 161474 3924 161480 3936
rect 110564 3896 161480 3924
rect 110564 3884 110570 3896
rect 161474 3884 161480 3896
rect 161532 3884 161538 3936
rect 25314 3816 25320 3868
rect 25372 3856 25378 3868
rect 59998 3856 60004 3868
rect 25372 3828 60004 3856
rect 25372 3816 25378 3828
rect 59998 3816 60004 3828
rect 60056 3816 60062 3868
rect 60826 3816 60832 3868
rect 60884 3856 60890 3868
rect 106366 3856 106372 3868
rect 60884 3828 106372 3856
rect 60884 3816 60890 3828
rect 106366 3816 106372 3828
rect 106424 3816 106430 3868
rect 106921 3859 106979 3865
rect 106921 3825 106933 3859
rect 106967 3856 106979 3859
rect 110414 3856 110420 3868
rect 106967 3828 110420 3856
rect 106967 3825 106979 3828
rect 106921 3819 106979 3825
rect 110414 3816 110420 3828
rect 110472 3816 110478 3868
rect 117041 3859 117099 3865
rect 117041 3825 117053 3859
rect 117087 3856 117099 3859
rect 160186 3856 160192 3868
rect 117087 3828 160192 3856
rect 117087 3825 117099 3828
rect 117041 3819 117099 3825
rect 160186 3816 160192 3828
rect 160244 3816 160250 3868
rect 8754 3748 8760 3800
rect 8812 3788 8818 3800
rect 25498 3788 25504 3800
rect 8812 3760 25504 3788
rect 8812 3748 8818 3760
rect 25498 3748 25504 3760
rect 25556 3748 25562 3800
rect 26510 3748 26516 3800
rect 26568 3788 26574 3800
rect 43438 3788 43444 3800
rect 26568 3760 43444 3788
rect 26568 3748 26574 3760
rect 43438 3748 43444 3760
rect 43496 3748 43502 3800
rect 45462 3748 45468 3800
rect 45520 3788 45526 3800
rect 83458 3788 83464 3800
rect 45520 3760 83464 3788
rect 45520 3748 45526 3760
rect 83458 3748 83464 3760
rect 83516 3748 83522 3800
rect 96246 3748 96252 3800
rect 96304 3788 96310 3800
rect 146294 3788 146300 3800
rect 96304 3760 146300 3788
rect 96304 3748 96310 3760
rect 146294 3748 146300 3760
rect 146352 3748 146358 3800
rect 2866 3680 2872 3732
rect 2924 3720 2930 3732
rect 15838 3720 15844 3732
rect 2924 3692 15844 3720
rect 2924 3680 2930 3692
rect 15838 3680 15844 3692
rect 15896 3680 15902 3732
rect 20622 3680 20628 3732
rect 20680 3720 20686 3732
rect 57238 3720 57244 3732
rect 20680 3692 57244 3720
rect 20680 3680 20686 3692
rect 57238 3680 57244 3692
rect 57296 3680 57302 3732
rect 67910 3680 67916 3732
rect 67968 3720 67974 3732
rect 67968 3692 108344 3720
rect 67968 3680 67974 3692
rect 15930 3612 15936 3664
rect 15988 3652 15994 3664
rect 55858 3652 55864 3664
rect 15988 3624 55864 3652
rect 15988 3612 15994 3624
rect 55858 3612 55864 3624
rect 55916 3612 55922 3664
rect 64322 3612 64328 3664
rect 64380 3652 64386 3664
rect 106921 3655 106979 3661
rect 106921 3652 106933 3655
rect 64380 3624 106933 3652
rect 64380 3612 64386 3624
rect 106921 3621 106933 3624
rect 106967 3621 106979 3655
rect 106921 3615 106979 3621
rect 7650 3544 7656 3596
rect 7708 3584 7714 3596
rect 8202 3584 8208 3596
rect 7708 3556 8208 3584
rect 7708 3544 7714 3556
rect 8202 3544 8208 3556
rect 8260 3544 8266 3596
rect 9950 3544 9956 3596
rect 10008 3584 10014 3596
rect 10962 3584 10968 3596
rect 10008 3556 10968 3584
rect 10008 3544 10014 3556
rect 10962 3544 10968 3556
rect 11020 3544 11026 3596
rect 11146 3544 11152 3596
rect 11204 3584 11210 3596
rect 52546 3584 52552 3596
rect 11204 3556 52552 3584
rect 11204 3544 11210 3556
rect 52546 3544 52552 3556
rect 52604 3544 52610 3596
rect 57238 3544 57244 3596
rect 57296 3584 57302 3596
rect 103514 3584 103520 3596
rect 57296 3556 103520 3584
rect 57296 3544 57302 3556
rect 103514 3544 103520 3556
rect 103572 3544 103578 3596
rect 108316 3584 108344 3692
rect 109310 3680 109316 3732
rect 109368 3720 109374 3732
rect 117041 3723 117099 3729
rect 117041 3720 117053 3723
rect 109368 3692 117053 3720
rect 109368 3680 109374 3692
rect 117041 3689 117053 3692
rect 117087 3689 117099 3723
rect 117041 3683 117099 3689
rect 117590 3680 117596 3732
rect 117648 3720 117654 3732
rect 169754 3720 169760 3732
rect 117648 3692 169760 3720
rect 117648 3680 117654 3692
rect 169754 3680 169760 3692
rect 169812 3680 169818 3732
rect 112806 3612 112812 3664
rect 112864 3652 112870 3664
rect 164234 3652 164240 3664
rect 112864 3624 164240 3652
rect 112864 3612 112870 3624
rect 164234 3612 164240 3624
rect 164292 3612 164298 3664
rect 114554 3584 114560 3596
rect 108316 3556 114560 3584
rect 114554 3544 114560 3556
rect 114612 3544 114618 3596
rect 116394 3544 116400 3596
rect 116452 3584 116458 3596
rect 168374 3584 168380 3596
rect 116452 3556 168380 3584
rect 116452 3544 116458 3556
rect 168374 3544 168380 3556
rect 168432 3544 168438 3596
rect 182082 3544 182088 3596
rect 182140 3584 182146 3596
rect 582190 3584 582196 3596
rect 182140 3556 582196 3584
rect 182140 3544 182146 3556
rect 582190 3544 582196 3556
rect 582248 3544 582254 3596
rect 6454 3476 6460 3528
rect 6512 3516 6518 3528
rect 47026 3516 47032 3528
rect 6512 3488 47032 3516
rect 6512 3476 6518 3488
rect 47026 3476 47032 3488
rect 47084 3476 47090 3528
rect 50154 3476 50160 3528
rect 50212 3516 50218 3528
rect 50982 3516 50988 3528
rect 50212 3488 50988 3516
rect 50212 3476 50218 3488
rect 50982 3476 50988 3488
rect 51040 3476 51046 3528
rect 53742 3476 53748 3528
rect 53800 3516 53806 3528
rect 95878 3516 95884 3528
rect 53800 3488 95884 3516
rect 53800 3476 53806 3488
rect 95878 3476 95884 3488
rect 95936 3476 95942 3528
rect 99834 3476 99840 3528
rect 99892 3516 99898 3528
rect 101398 3516 101404 3528
rect 99892 3488 101404 3516
rect 99892 3476 99898 3488
rect 101398 3476 101404 3488
rect 101456 3476 101462 3528
rect 103330 3476 103336 3528
rect 103388 3516 103394 3528
rect 154574 3516 154580 3528
rect 103388 3488 154580 3516
rect 103388 3476 103394 3488
rect 154574 3476 154580 3488
rect 154632 3476 154638 3528
rect 183462 3476 183468 3528
rect 183520 3516 183526 3528
rect 583386 3516 583392 3528
rect 183520 3488 583392 3516
rect 183520 3476 183526 3488
rect 583386 3476 583392 3488
rect 583444 3476 583450 3528
rect 5258 3408 5264 3460
rect 5316 3448 5322 3460
rect 45554 3448 45560 3460
rect 5316 3420 45560 3448
rect 5316 3408 5322 3420
rect 45554 3408 45560 3420
rect 45612 3408 45618 3460
rect 52546 3408 52552 3460
rect 52604 3448 52610 3460
rect 66898 3448 66904 3460
rect 52604 3420 66904 3448
rect 52604 3408 52610 3420
rect 66898 3408 66904 3420
rect 66956 3408 66962 3460
rect 69106 3408 69112 3460
rect 69164 3448 69170 3460
rect 70302 3448 70308 3460
rect 69164 3420 70308 3448
rect 69164 3408 69170 3420
rect 70302 3408 70308 3420
rect 70360 3408 70366 3460
rect 71498 3408 71504 3460
rect 71556 3448 71562 3460
rect 71556 3420 103514 3448
rect 71556 3408 71562 3420
rect 566 3340 572 3392
rect 624 3380 630 3392
rect 2038 3380 2044 3392
rect 624 3352 2044 3380
rect 624 3340 630 3352
rect 2038 3340 2044 3352
rect 2096 3340 2102 3392
rect 18230 3340 18236 3392
rect 18288 3380 18294 3392
rect 21450 3380 21456 3392
rect 18288 3352 21456 3380
rect 18288 3340 18294 3352
rect 21450 3340 21456 3352
rect 21508 3340 21514 3392
rect 24210 3340 24216 3392
rect 24268 3380 24274 3392
rect 24762 3380 24768 3392
rect 24268 3352 24768 3380
rect 24268 3340 24274 3352
rect 24762 3340 24768 3352
rect 24820 3340 24826 3392
rect 32398 3340 32404 3392
rect 32456 3380 32462 3392
rect 33042 3380 33048 3392
rect 32456 3352 33048 3380
rect 32456 3340 32462 3352
rect 33042 3340 33048 3352
rect 33100 3340 33106 3392
rect 35986 3340 35992 3392
rect 36044 3380 36050 3392
rect 37182 3380 37188 3392
rect 36044 3352 37188 3380
rect 36044 3340 36050 3352
rect 37182 3340 37188 3352
rect 37240 3340 37246 3392
rect 41874 3340 41880 3392
rect 41932 3380 41938 3392
rect 42702 3380 42708 3392
rect 41932 3352 42708 3380
rect 41932 3340 41938 3352
rect 42702 3340 42708 3352
rect 42760 3340 42766 3392
rect 66714 3340 66720 3392
rect 66772 3380 66778 3392
rect 75178 3380 75184 3392
rect 66772 3352 75184 3380
rect 66772 3340 66778 3352
rect 75178 3340 75184 3352
rect 75236 3340 75242 3392
rect 84470 3340 84476 3392
rect 84528 3380 84534 3392
rect 86218 3380 86224 3392
rect 84528 3352 86224 3380
rect 84528 3340 84534 3352
rect 86218 3340 86224 3352
rect 86276 3340 86282 3392
rect 103486 3380 103514 3420
rect 106918 3408 106924 3460
rect 106976 3448 106982 3460
rect 108298 3448 108304 3460
rect 106976 3420 108304 3448
rect 106976 3408 106982 3420
rect 108298 3408 108304 3420
rect 108356 3408 108362 3460
rect 114002 3408 114008 3460
rect 114060 3448 114066 3460
rect 114462 3448 114468 3460
rect 114060 3420 114468 3448
rect 114060 3408 114066 3420
rect 114462 3408 114468 3420
rect 114520 3408 114526 3460
rect 115198 3408 115204 3460
rect 115256 3448 115262 3460
rect 115842 3448 115848 3460
rect 115256 3420 115848 3448
rect 115256 3408 115262 3420
rect 115842 3408 115848 3420
rect 115900 3408 115906 3460
rect 121086 3408 121092 3460
rect 121144 3448 121150 3460
rect 173894 3448 173900 3460
rect 121144 3420 173900 3448
rect 121144 3408 121150 3420
rect 173894 3408 173900 3420
rect 173952 3408 173958 3460
rect 180702 3408 180708 3460
rect 180760 3448 180766 3460
rect 580994 3448 581000 3460
rect 180760 3420 581000 3448
rect 180760 3408 180766 3420
rect 580994 3408 581000 3420
rect 581052 3408 581058 3460
rect 118878 3380 118884 3392
rect 103486 3352 118884 3380
rect 118878 3340 118884 3352
rect 118936 3340 118942 3392
rect 1670 3272 1676 3324
rect 1728 3312 1734 3324
rect 6178 3312 6184 3324
rect 1728 3284 6184 3312
rect 1728 3272 1734 3284
rect 6178 3272 6184 3284
rect 6236 3272 6242 3324
rect 33594 3272 33600 3324
rect 33652 3312 33658 3324
rect 40126 3312 40132 3324
rect 33652 3284 40132 3312
rect 33652 3272 33658 3284
rect 40126 3272 40132 3284
rect 40184 3272 40190 3324
rect 44266 3272 44272 3324
rect 44324 3312 44330 3324
rect 51074 3312 51080 3324
rect 44324 3284 51080 3312
rect 44324 3272 44330 3284
rect 51074 3272 51080 3284
rect 51132 3272 51138 3324
rect 65518 3272 65524 3324
rect 65576 3312 65582 3324
rect 66162 3312 66168 3324
rect 65576 3284 66168 3312
rect 65576 3272 65582 3284
rect 66162 3272 66168 3284
rect 66220 3272 66226 3324
rect 58434 3136 58440 3188
rect 58492 3176 58498 3188
rect 61930 3176 61936 3188
rect 58492 3148 61936 3176
rect 58492 3136 58498 3148
rect 61930 3136 61936 3148
rect 61988 3136 61994 3188
rect 85666 3136 85672 3188
rect 85724 3176 85730 3188
rect 90266 3176 90272 3188
rect 85724 3148 90272 3176
rect 85724 3136 85730 3148
rect 90266 3136 90272 3148
rect 90324 3136 90330 3188
rect 17034 3068 17040 3120
rect 17092 3108 17098 3120
rect 19978 3108 19984 3120
rect 17092 3080 19984 3108
rect 17092 3068 17098 3080
rect 19978 3068 19984 3080
rect 20036 3068 20042 3120
rect 46658 2932 46664 2984
rect 46716 2972 46722 2984
rect 54478 2972 54484 2984
rect 46716 2944 54484 2972
rect 46716 2932 46722 2944
rect 54478 2932 54484 2944
rect 54536 2932 54542 2984
rect 87966 2932 87972 2984
rect 88024 2972 88030 2984
rect 88426 2972 88432 2984
rect 88024 2944 88432 2972
rect 88024 2932 88030 2944
rect 88426 2932 88432 2944
rect 88484 2932 88490 2984
rect 12342 2864 12348 2916
rect 12400 2904 12406 2916
rect 17218 2904 17224 2916
rect 12400 2876 17224 2904
rect 12400 2864 12406 2876
rect 17218 2864 17224 2876
rect 17276 2864 17282 2916
rect 124674 2796 124680 2848
rect 124732 2836 124738 2848
rect 128538 2836 128544 2848
rect 124732 2808 128544 2836
rect 124732 2796 124738 2808
rect 128538 2796 128544 2808
rect 128596 2796 128602 2848
<< via1 >>
rect 201500 702992 201552 703044
rect 202788 702992 202840 703044
rect 229744 700952 229796 701004
rect 267648 700952 267700 701004
rect 211804 700884 211856 700936
rect 332508 700884 332560 700936
rect 220084 700816 220136 700868
rect 348792 700816 348844 700868
rect 193864 700748 193916 700800
rect 364984 700748 365036 700800
rect 209044 700680 209096 700732
rect 397460 700680 397512 700732
rect 215944 700612 215996 700664
rect 413652 700612 413704 700664
rect 191104 700544 191156 700596
rect 429844 700544 429896 700596
rect 204904 700476 204956 700528
rect 462320 700476 462372 700528
rect 170312 700408 170364 700460
rect 176844 700408 176896 700460
rect 198004 700408 198056 700460
rect 235172 700408 235224 700460
rect 238024 700408 238076 700460
rect 527180 700408 527232 700460
rect 137836 700340 137888 700392
rect 176752 700340 176804 700392
rect 189724 700340 189776 700392
rect 494796 700340 494848 700392
rect 89168 700272 89220 700324
rect 176660 700272 176712 700324
rect 185584 700272 185636 700324
rect 559656 700272 559708 700324
rect 24308 699660 24360 699712
rect 24768 699660 24820 699712
rect 39856 699660 39908 699712
rect 40500 699660 40552 699712
rect 71780 699660 71832 699712
rect 72976 699660 73028 699712
rect 105452 699660 105504 699712
rect 106188 699660 106240 699712
rect 196624 696940 196676 696992
rect 580172 696940 580224 696992
rect 2780 683612 2832 683664
rect 6184 683612 6236 683664
rect 182824 670692 182876 670744
rect 580172 670692 580224 670744
rect 3516 656888 3568 656940
rect 21364 656888 21416 656940
rect 200764 643084 200816 643136
rect 580172 643084 580224 643136
rect 3516 632068 3568 632120
rect 15844 632068 15896 632120
rect 214564 630640 214616 630692
rect 579988 630640 580040 630692
rect 180064 616836 180116 616888
rect 580172 616836 580224 616888
rect 3332 605820 3384 605872
rect 25504 605820 25556 605872
rect 226984 590656 227036 590708
rect 580172 590656 580224 590708
rect 3332 579640 3384 579692
rect 10324 579640 10376 579692
rect 231124 563048 231176 563100
rect 579896 563048 579948 563100
rect 3332 553392 3384 553444
rect 28264 553392 28316 553444
rect 269764 536800 269816 536852
rect 580172 536800 580224 536852
rect 3332 527144 3384 527196
rect 13084 527144 13136 527196
rect 267004 524424 267056 524476
rect 580172 524424 580224 524476
rect 3332 514768 3384 514820
rect 35164 514768 35216 514820
rect 265624 510620 265676 510672
rect 580172 510620 580224 510672
rect 2872 500964 2924 501016
rect 31024 500964 31076 501016
rect 268384 484372 268436 484424
rect 580172 484372 580224 484424
rect 3332 474716 3384 474768
rect 14464 474716 14516 474768
rect 153200 472608 153252 472660
rect 176936 472608 176988 472660
rect 3332 462340 3384 462392
rect 19984 462340 20036 462392
rect 479524 456764 479576 456816
rect 579620 456764 579672 456816
rect 3332 448536 3384 448588
rect 32404 448536 32456 448588
rect 39764 425688 39816 425740
rect 71780 425688 71832 425740
rect 106188 425688 106240 425740
rect 177028 425688 177080 425740
rect 3148 422288 3200 422340
rect 17224 422288 17276 422340
rect 486424 418140 486476 418192
rect 579712 418140 579764 418192
rect 482284 404336 482336 404388
rect 580172 404336 580224 404388
rect 3332 397468 3384 397520
rect 33784 397468 33836 397520
rect 483664 378156 483716 378208
rect 580172 378156 580224 378208
rect 294604 376728 294656 376780
rect 337660 376728 337712 376780
rect 262864 375368 262916 375420
rect 337752 375368 337804 375420
rect 291844 372580 291896 372632
rect 337476 372580 337528 372632
rect 3332 371220 3384 371272
rect 20076 371220 20128 371272
rect 261484 369928 261536 369980
rect 337476 369928 337528 369980
rect 35624 369860 35676 369912
rect 37924 369860 37976 369912
rect 258724 369860 258776 369912
rect 337752 369860 337804 369912
rect 195888 367072 195940 367124
rect 337476 367072 337528 367124
rect 485044 364352 485096 364404
rect 580172 364352 580224 364404
rect 480904 351908 480956 351960
rect 580172 351908 580224 351960
rect 187608 349120 187660 349172
rect 337752 349120 337804 349172
rect 35808 347828 35860 347880
rect 37648 347828 37700 347880
rect 254584 347760 254636 347812
rect 337660 347760 337712 347812
rect 3056 345040 3108 345092
rect 35256 345040 35308 345092
rect 35164 339396 35216 339448
rect 146300 339396 146352 339448
rect 3424 339328 3476 339380
rect 133880 339328 133932 339380
rect 3516 339260 3568 339312
rect 138020 339260 138072 339312
rect 100668 339192 100720 339244
rect 238024 339192 238076 339244
rect 3608 339124 3660 339176
rect 142160 339124 142212 339176
rect 3792 339056 3844 339108
rect 157340 339056 157392 339108
rect 38752 338988 38804 339040
rect 202972 338988 203024 339040
rect 38384 338920 38436 338972
rect 240692 338920 240744 338972
rect 97908 338852 97960 338904
rect 580264 338852 580316 338904
rect 89536 338784 89588 338836
rect 580356 338784 580408 338836
rect 82728 338716 82780 338768
rect 580540 338716 580592 338768
rect 39856 338648 39908 338700
rect 128360 338648 128412 338700
rect 121368 338580 121420 338632
rect 176844 338580 176896 338632
rect 38568 338036 38620 338088
rect 337384 338036 337436 338088
rect 42064 337832 42116 337884
rect 379520 337832 379572 337884
rect 50344 337764 50396 337816
rect 394700 337764 394752 337816
rect 78588 337696 78640 337748
rect 56508 337628 56560 337680
rect 61384 337628 61436 337680
rect 77208 337628 77260 337680
rect 79324 337628 79376 337680
rect 122748 337696 122800 337748
rect 176752 337696 176804 337748
rect 388444 337696 388496 337748
rect 391940 337696 391992 337748
rect 126244 337628 126296 337680
rect 143448 337628 143500 337680
rect 241520 337628 241572 337680
rect 367744 337628 367796 337680
rect 369860 337628 369912 337680
rect 387064 337628 387116 337680
rect 389180 337628 389232 337680
rect 118608 337560 118660 337612
rect 237748 337560 237800 337612
rect 117228 337492 117280 337544
rect 237656 337492 237708 337544
rect 355324 337492 355376 337544
rect 372620 337492 372672 337544
rect 104808 337424 104860 337476
rect 237564 337424 237616 337476
rect 364984 337424 365036 337476
rect 397460 337424 397512 337476
rect 43444 337356 43496 337408
rect 96620 337356 96672 337408
rect 99288 337356 99340 337408
rect 236644 337356 236696 337408
rect 349804 337356 349856 337408
rect 385040 337356 385092 337408
rect 93584 337288 93636 337340
rect 232504 337288 232556 337340
rect 352564 337288 352616 337340
rect 387800 337356 387852 337408
rect 385684 337288 385736 337340
rect 390560 337288 390612 337340
rect 89628 337220 89680 337272
rect 238300 337220 238352 337272
rect 287704 337220 287756 337272
rect 382280 337220 382332 337272
rect 84016 337152 84068 337204
rect 238208 337152 238260 337204
rect 255964 337152 256016 337204
rect 371240 337152 371292 337204
rect 382924 337152 382976 337204
rect 386420 337152 386472 337204
rect 40500 337084 40552 337136
rect 60740 337084 60792 337136
rect 67548 337084 67600 337136
rect 236736 337084 236788 337136
rect 249064 337084 249116 337136
rect 375380 337084 375432 337136
rect 381544 337084 381596 337136
rect 386512 337084 386564 337136
rect 38384 337016 38436 337068
rect 59360 337016 59412 337068
rect 66168 337016 66220 337068
rect 239404 337016 239456 337068
rect 251824 337016 251876 337068
rect 433340 337016 433392 337068
rect 46204 336948 46256 337000
rect 379428 336948 379480 337000
rect 379520 336948 379572 337000
rect 387800 336948 387852 337000
rect 411904 336948 411956 337000
rect 440240 336948 440292 337000
rect 48964 336880 49016 336932
rect 383752 336880 383804 336932
rect 402244 336880 402296 336932
rect 407120 336880 407172 336932
rect 409144 336880 409196 336932
rect 425060 336880 425112 336932
rect 384948 336812 385000 336864
rect 396080 336812 396132 336864
rect 399484 336812 399536 336864
rect 405740 336812 405792 336864
rect 406384 336812 406436 336864
rect 422944 336812 422996 336864
rect 40316 336744 40368 336796
rect 57980 336744 58032 336796
rect 70308 336744 70360 336796
rect 75184 336744 75236 336796
rect 95148 336744 95200 336796
rect 106924 336744 106976 336796
rect 351184 336744 351236 336796
rect 364524 336744 364576 336796
rect 373264 336744 373316 336796
rect 378140 336744 378192 336796
rect 391204 336744 391256 336796
rect 393320 336744 393372 336796
rect 290464 336608 290516 336660
rect 390560 336608 390612 336660
rect 81348 336540 81400 336592
rect 173164 336540 173216 336592
rect 250444 336540 250496 336592
rect 376852 336540 376904 336592
rect 131028 336472 131080 336524
rect 225604 336472 225656 336524
rect 234528 336472 234580 336524
rect 384948 336472 385000 336524
rect 129648 336404 129700 336456
rect 175924 336404 175976 336456
rect 223488 336404 223540 336456
rect 379520 336404 379572 336456
rect 81256 336336 81308 336388
rect 177304 336336 177356 336388
rect 243544 336336 243596 336388
rect 403256 336336 403308 336388
rect 37096 336268 37148 336320
rect 98000 336268 98052 336320
rect 121276 336268 121328 336320
rect 220820 336268 220872 336320
rect 244924 336268 244976 336320
rect 409880 336268 409932 336320
rect 37188 336200 37240 336252
rect 75920 336200 75972 336252
rect 96528 336200 96580 336252
rect 207664 336200 207716 336252
rect 213828 336200 213880 336252
rect 397460 336200 397512 336252
rect 19984 336132 20036 336184
rect 150440 336132 150492 336184
rect 247684 336132 247736 336184
rect 443000 336132 443052 336184
rect 35716 336064 35768 336116
rect 371240 336064 371292 336116
rect 38752 335996 38804 336048
rect 382372 335996 382424 336048
rect 82176 334568 82228 334620
rect 178684 334568 178736 334620
rect 71320 331848 71372 331900
rect 238760 331848 238812 331900
rect 68744 324300 68796 324352
rect 579988 324300 580040 324352
rect 3424 318792 3476 318844
rect 158720 318792 158772 318844
rect 70308 311856 70360 311908
rect 580172 311856 580224 311908
rect 3424 304988 3476 305040
rect 161480 304988 161532 305040
rect 67548 298120 67600 298172
rect 580172 298120 580224 298172
rect 3424 292544 3476 292596
rect 160100 292544 160152 292596
rect 66168 271872 66220 271924
rect 580172 271872 580224 271924
rect 216588 269764 216640 269816
rect 399576 269764 399628 269816
rect 10324 268404 10376 268456
rect 139400 268404 139452 268456
rect 20076 268336 20128 268388
rect 154580 268336 154632 268388
rect 108856 266976 108908 267028
rect 215944 266976 215996 267028
rect 3056 266364 3108 266416
rect 162860 266364 162912 266416
rect 32404 262896 32456 262948
rect 149060 262896 149112 262948
rect 38844 262828 38896 262880
rect 195980 262828 196032 262880
rect 66076 258068 66128 258120
rect 580172 258068 580224 258120
rect 3424 253920 3476 253972
rect 165620 253920 165672 253972
rect 86776 253172 86828 253224
rect 231124 253172 231176 253224
rect 91008 252152 91060 252204
rect 204996 252152 205048 252204
rect 106924 252084 106976 252136
rect 229100 252084 229152 252136
rect 85488 252016 85540 252068
rect 219440 252016 219492 252068
rect 79324 251948 79376 252000
rect 213920 251948 213972 252000
rect 64788 251880 64840 251932
rect 237932 251880 237984 251932
rect 35348 251812 35400 251864
rect 393412 251812 393464 251864
rect 25504 250860 25556 250912
rect 136640 250860 136692 250912
rect 119804 250792 119856 250844
rect 282920 250792 282972 250844
rect 84292 250724 84344 250776
rect 267004 250724 267056 250776
rect 35532 250656 35584 250708
rect 369952 250656 370004 250708
rect 77300 250588 77352 250640
rect 486424 250588 486476 250640
rect 71780 250520 71832 250572
rect 483664 250520 483716 250572
rect 99380 250452 99432 250504
rect 542360 250452 542412 250504
rect 117320 249704 117372 249756
rect 201500 249704 201552 249756
rect 36636 249636 36688 249688
rect 122840 249636 122892 249688
rect 100760 249568 100812 249620
rect 189724 249568 189776 249620
rect 110420 249500 110472 249552
rect 211804 249500 211856 249552
rect 95240 249432 95292 249484
rect 196624 249432 196676 249484
rect 106280 249364 106332 249416
rect 209044 249364 209096 249416
rect 102140 249296 102192 249348
rect 204904 249296 204956 249348
rect 114560 249228 114612 249280
rect 229744 249228 229796 249280
rect 86960 249160 87012 249212
rect 226984 249160 227036 249212
rect 82820 249092 82872 249144
rect 269764 249092 269816 249144
rect 35440 249024 35492 249076
rect 380992 249024 381044 249076
rect 105728 248344 105780 248396
rect 191104 248344 191156 248396
rect 98092 248276 98144 248328
rect 185584 248276 185636 248328
rect 90364 248208 90416 248260
rect 180064 248208 180116 248260
rect 91652 248140 91704 248192
rect 200764 248140 200816 248192
rect 6184 248072 6236 248124
rect 132592 248072 132644 248124
rect 86868 248004 86920 248056
rect 241704 248004 241756 248056
rect 82636 247936 82688 247988
rect 265624 247936 265676 247988
rect 80152 247868 80204 247920
rect 268384 247868 268436 247920
rect 78864 247800 78916 247852
rect 479524 247800 479576 247852
rect 75092 247732 75144 247784
rect 482284 247732 482336 247784
rect 71228 247664 71280 247716
rect 480904 247664 480956 247716
rect 109592 247596 109644 247648
rect 193864 247596 193916 247648
rect 36820 247528 36872 247580
rect 113180 247528 113232 247580
rect 94228 246848 94280 246900
rect 182824 246848 182876 246900
rect 24768 246780 24820 246832
rect 131304 246780 131356 246832
rect 93676 246712 93728 246764
rect 208032 246712 208084 246764
rect 108948 246644 109000 246696
rect 239312 246644 239364 246696
rect 60648 246576 60700 246628
rect 192668 246576 192720 246628
rect 57888 246508 57940 246560
rect 191380 246508 191432 246560
rect 38200 246440 38252 246492
rect 186320 246440 186372 246492
rect 3700 246372 3752 246424
rect 154304 246372 154356 246424
rect 38660 246304 38712 246356
rect 199108 246304 199160 246356
rect 21364 245556 21416 245608
rect 133880 245556 133932 245608
rect 31024 245488 31076 245540
rect 145380 245488 145432 245540
rect 146208 245488 146260 245540
rect 241612 245488 241664 245540
rect 33784 245420 33836 245472
rect 153016 245420 153068 245472
rect 92940 245352 92992 245404
rect 214564 245352 214616 245404
rect 102048 245284 102100 245336
rect 239220 245284 239272 245336
rect 35256 245216 35308 245268
rect 156880 245216 156932 245268
rect 205456 245216 205508 245268
rect 349804 245216 349856 245268
rect 68836 245148 68888 245200
rect 238944 245148 238996 245200
rect 8208 245080 8260 245132
rect 130016 245080 130068 245132
rect 231032 245080 231084 245132
rect 437480 245080 437532 245132
rect 39580 245012 39632 245064
rect 89720 245012 89772 245064
rect 104440 245012 104492 245064
rect 477500 245012 477552 245064
rect 73804 244944 73856 244996
rect 485044 244944 485096 244996
rect 76380 244876 76432 244928
rect 580448 244876 580500 244928
rect 28264 244808 28316 244860
rect 141516 244808 141568 244860
rect 36912 244740 36964 244792
rect 104900 244740 104952 244792
rect 112168 244740 112220 244792
rect 220084 244740 220136 244792
rect 119988 244672 120040 244724
rect 218060 244672 218112 244724
rect 117228 243924 117280 243976
rect 198004 243924 198056 243976
rect 198096 243924 198148 243976
rect 249064 243924 249116 243976
rect 15844 243856 15896 243908
rect 136456 243856 136508 243908
rect 142068 243856 142120 243908
rect 240600 243856 240652 243908
rect 13084 243788 13136 243840
rect 144092 243788 144144 243840
rect 193956 243788 194008 243840
rect 355324 243788 355376 243840
rect 113456 243720 113508 243772
rect 299480 243720 299532 243772
rect 14464 243652 14516 243704
rect 147956 243652 148008 243704
rect 225972 243652 226024 243704
rect 430580 243652 430632 243704
rect 17224 243584 17276 243636
rect 151820 243584 151872 243636
rect 236184 243584 236236 243636
rect 445760 243584 445812 243636
rect 85488 243516 85540 243568
rect 579620 243516 579672 243568
rect 15936 243448 15988 243500
rect 167092 243448 167144 243500
rect 28264 243380 28316 243432
rect 179880 243380 179932 243432
rect 17316 243312 17368 243364
rect 170956 243312 171008 243364
rect 19984 243244 20036 243296
rect 174820 243244 174872 243296
rect 21364 243176 21416 243228
rect 182456 243176 182508 243228
rect 6184 243108 6236 243160
rect 178592 243108 178644 243160
rect 48228 243040 48280 243092
rect 268384 243040 268436 243092
rect 44364 242972 44416 243024
rect 267004 242972 267056 243024
rect 41788 242904 41840 242956
rect 273904 242904 273956 242956
rect 81440 242836 81492 242888
rect 82728 242836 82780 242888
rect 82820 242836 82872 242888
rect 84016 242836 84068 242888
rect 84292 242836 84344 242888
rect 85304 242836 85356 242888
rect 86960 242836 87012 242888
rect 87880 242836 87932 242888
rect 96804 242836 96856 242888
rect 97908 242836 97960 242888
rect 99380 242836 99432 242888
rect 100300 242836 100352 242888
rect 100760 242836 100812 242888
rect 101956 242836 102008 242888
rect 102140 242836 102192 242888
rect 103152 242836 103204 242888
rect 106280 242836 106332 242888
rect 107016 242836 107068 242888
rect 117320 242836 117372 242888
rect 118516 242836 118568 242888
rect 126244 242836 126296 242888
rect 240508 242836 240560 242888
rect 79968 242768 80020 242820
rect 96344 242700 96396 242752
rect 232320 242700 232372 242752
rect 233608 242768 233660 242820
rect 234528 242768 234580 242820
rect 238116 242768 238168 242820
rect 237472 242700 237524 242752
rect 398104 242700 398156 242752
rect 99380 242632 99432 242684
rect 100668 242632 100720 242684
rect 115940 242632 115992 242684
rect 119804 242632 119856 242684
rect 177304 242632 177356 242684
rect 215668 242632 215720 242684
rect 216588 242632 216640 242684
rect 220820 242632 220872 242684
rect 175924 242564 175976 242616
rect 224684 242564 224736 242616
rect 225604 242632 225656 242684
rect 227168 242632 227220 242684
rect 382924 242632 382976 242684
rect 228456 242564 228508 242616
rect 391204 242564 391256 242616
rect 64880 242496 64932 242548
rect 66168 242496 66220 242548
rect 124956 242496 125008 242548
rect 177028 242496 177080 242548
rect 204996 242496 205048 242548
rect 206744 242496 206796 242548
rect 207664 242496 207716 242548
rect 210608 242496 210660 242548
rect 211896 242496 211948 242548
rect 375472 242496 375524 242548
rect 75184 242428 75236 242480
rect 202880 242428 202932 242480
rect 209320 242428 209372 242480
rect 374000 242428 374052 242480
rect 39764 242360 39816 242412
rect 126244 242360 126296 242412
rect 200396 242360 200448 242412
rect 366364 242360 366416 242412
rect 63592 242292 63644 242344
rect 85488 242292 85540 242344
rect 123668 242292 123720 242344
rect 176936 242292 176988 242344
rect 190092 242292 190144 242344
rect 356060 242292 356112 242344
rect 36544 242224 36596 242276
rect 125600 242224 125652 242276
rect 127440 242224 127492 242276
rect 176660 242224 176712 242276
rect 188896 242224 188948 242276
rect 363052 242224 363104 242276
rect 35256 242156 35308 242208
rect 376760 242156 376812 242208
rect 133788 242088 133840 242140
rect 239496 242088 239548 242140
rect 136548 242020 136600 242072
rect 240140 242020 240192 242072
rect 61016 241952 61068 242004
rect 96528 241952 96580 242004
rect 178684 241952 178736 242004
rect 218244 241952 218296 242004
rect 234896 241952 234948 242004
rect 247684 241952 247736 242004
rect 53288 241884 53340 241936
rect 128820 241884 128872 241936
rect 173164 241884 173216 241936
rect 201592 241884 201644 241936
rect 216956 241884 217008 241936
rect 62304 241816 62356 241868
rect 178040 241816 178092 241868
rect 58440 241748 58492 241800
rect 177396 241748 177448 241800
rect 46940 241680 46992 241732
rect 175188 241680 175240 241732
rect 3424 241612 3476 241664
rect 164516 241612 164568 241664
rect 13084 241544 13136 241596
rect 181168 241544 181220 241596
rect 14464 241476 14516 241528
rect 185032 241476 185084 241528
rect 38568 241408 38620 241460
rect 39304 241408 39356 241460
rect 39396 241408 39448 241460
rect 74632 241408 74684 241460
rect 39120 241340 39172 241392
rect 85672 241340 85724 241392
rect 39212 241272 39264 241324
rect 87052 241272 87104 241324
rect 99104 241272 99156 241324
rect 238852 241272 238904 241324
rect 39488 241204 39540 241256
rect 91192 241204 91244 241256
rect 92388 241204 92440 241256
rect 238024 241204 238076 241256
rect 68928 241136 68980 241188
rect 239128 241136 239180 241188
rect 38844 241068 38896 241120
rect 365720 241068 365772 241120
rect 37004 241000 37056 241052
rect 367192 241000 367244 241052
rect 38108 240932 38160 240984
rect 368480 240932 368532 240984
rect 37740 240864 37792 240916
rect 381544 240864 381596 240916
rect 36728 240796 36780 240848
rect 412640 240796 412692 240848
rect 61384 240728 61436 240780
rect 240416 240728 240468 240780
rect 39028 240116 39080 240168
rect 39396 240116 39448 240168
rect 168472 240048 168524 240100
rect 580172 240048 580224 240100
rect 38016 239980 38068 240032
rect 42064 239980 42116 240032
rect 236644 239980 236696 240032
rect 237840 239980 237892 240032
rect 240876 239980 240928 240032
rect 37924 239912 37976 239964
rect 46204 239912 46256 239964
rect 171876 239955 171928 239964
rect 37832 239844 37884 239896
rect 48964 239844 49016 239896
rect 33784 239776 33836 239828
rect 39396 239708 39448 239760
rect 39580 239708 39632 239760
rect 40132 239708 40184 239760
rect 43444 239708 43496 239760
rect 50344 239844 50396 239896
rect 171876 239921 171885 239955
rect 171885 239921 171919 239955
rect 171919 239921 171928 239955
rect 171876 239912 171928 239921
rect 236736 239912 236788 239964
rect 240324 239912 240376 239964
rect 139308 239844 139360 239896
rect 239036 239844 239088 239896
rect 183560 239776 183612 239828
rect 232504 239776 232556 239828
rect 49608 239751 49660 239760
rect 49608 239717 49617 239751
rect 49617 239717 49651 239751
rect 49651 239717 49660 239751
rect 49608 239708 49660 239717
rect 52368 239751 52420 239760
rect 52368 239717 52377 239751
rect 52377 239717 52411 239751
rect 52411 239717 52420 239751
rect 52368 239708 52420 239717
rect 54852 239751 54904 239760
rect 54852 239717 54861 239751
rect 54861 239717 54895 239751
rect 54895 239717 54904 239751
rect 54852 239708 54904 239717
rect 56232 239751 56284 239760
rect 56232 239717 56241 239751
rect 56241 239717 56275 239751
rect 56275 239717 56284 239751
rect 56232 239708 56284 239717
rect 57520 239751 57572 239760
rect 57520 239717 57529 239751
rect 57529 239717 57563 239751
rect 57563 239717 57572 239751
rect 57520 239708 57572 239717
rect 57704 239751 57756 239760
rect 57704 239717 57713 239751
rect 57713 239717 57747 239751
rect 57747 239717 57756 239751
rect 57704 239708 57756 239717
rect 59176 239751 59228 239760
rect 59176 239717 59185 239751
rect 59185 239717 59219 239751
rect 59219 239717 59228 239751
rect 59176 239708 59228 239717
rect 60096 239751 60148 239760
rect 60096 239717 60105 239751
rect 60105 239717 60139 239751
rect 60139 239717 60148 239751
rect 60096 239708 60148 239717
rect 62120 239751 62172 239760
rect 62120 239717 62129 239751
rect 62129 239717 62163 239751
rect 62163 239717 62172 239751
rect 62120 239708 62172 239717
rect 73436 239751 73488 239760
rect 73436 239717 73445 239751
rect 73445 239717 73479 239751
rect 73479 239717 73488 239751
rect 73436 239708 73488 239717
rect 75828 239751 75880 239760
rect 75828 239717 75837 239751
rect 75837 239717 75871 239751
rect 75871 239717 75880 239751
rect 75828 239708 75880 239717
rect 82912 239751 82964 239760
rect 82912 239717 82921 239751
rect 82921 239717 82955 239751
rect 82955 239717 82964 239751
rect 82912 239708 82964 239717
rect 96528 239708 96580 239760
rect 128820 239751 128872 239760
rect 128820 239717 128829 239751
rect 128829 239717 128863 239751
rect 128863 239717 128872 239751
rect 128820 239708 128872 239717
rect 31024 239640 31076 239692
rect 173164 239708 173216 239760
rect 175188 239708 175240 239760
rect 168472 239683 168524 239692
rect 168472 239649 168481 239683
rect 168481 239649 168515 239683
rect 168515 239649 168524 239683
rect 168472 239640 168524 239649
rect 169300 239683 169352 239692
rect 169300 239649 169309 239683
rect 169309 239649 169343 239683
rect 169343 239649 169352 239683
rect 169300 239640 169352 239649
rect 25504 239572 25556 239624
rect 175740 239640 175792 239692
rect 178040 239708 178092 239760
rect 580632 239708 580684 239760
rect 177028 239683 177080 239692
rect 177028 239649 177037 239683
rect 177037 239649 177071 239683
rect 177071 239649 177080 239683
rect 177028 239640 177080 239649
rect 177396 239640 177448 239692
rect 580540 239640 580592 239692
rect 24124 239504 24176 239556
rect 580264 239504 580316 239556
rect 40224 239436 40276 239488
rect 580448 239436 580500 239488
rect 38936 239368 38988 239420
rect 580356 239368 580408 239420
rect 10324 239300 10376 239352
rect 7564 239232 7616 239284
rect 3424 239164 3476 239216
rect 38660 239096 38712 239148
rect 272524 239096 272576 239148
rect 269764 239028 269816 239080
rect 280804 238960 280856 239012
rect 279424 238892 279476 238944
rect 284944 238824 284996 238876
rect 341524 238756 341576 238808
rect 38568 238688 38620 238740
rect 40224 238688 40276 238740
rect 241152 238688 241204 238740
rect 364984 238688 365036 238740
rect 38292 238144 38344 238196
rect 357440 238144 357492 238196
rect 580356 235492 580408 235544
rect 580724 235492 580776 235544
rect 38200 232772 38252 232824
rect 40408 232772 40460 232824
rect 38292 231956 38344 232008
rect 38568 231956 38620 232008
rect 238300 229032 238352 229084
rect 240600 229032 240652 229084
rect 240232 226992 240284 227044
rect 240416 226992 240468 227044
rect 240324 226040 240376 226092
rect 240324 225836 240376 225888
rect 239404 224748 239456 224800
rect 240416 224748 240468 224800
rect 3332 215228 3384 215280
rect 15936 215228 15988 215280
rect 241244 213868 241296 213920
rect 251824 213868 251876 213920
rect 241428 208292 241480 208344
rect 388444 208292 388496 208344
rect 272524 206932 272576 206984
rect 579804 206932 579856 206984
rect 285680 204892 285732 204944
rect 427820 204892 427872 204944
rect 3056 202784 3108 202836
rect 10324 202784 10376 202836
rect 241428 202784 241480 202836
rect 285680 202784 285732 202836
rect 241428 198636 241480 198688
rect 387064 198636 387116 198688
rect 238208 195916 238260 195968
rect 240140 195916 240192 195968
rect 280804 193128 280856 193180
rect 579620 193128 579672 193180
rect 3516 188844 3568 188896
rect 7564 188844 7616 188896
rect 241428 187620 241480 187672
rect 417424 187620 417476 187672
rect 285680 185580 285732 185632
rect 415400 185580 415452 185632
rect 241428 183472 241480 183524
rect 285680 183472 285732 183524
rect 241244 173612 241296 173664
rect 244924 173612 244976 173664
rect 35624 169464 35676 169516
rect 37832 169464 37884 169516
rect 269764 166948 269816 167000
rect 580172 166948 580224 167000
rect 3240 164160 3292 164212
rect 17316 164160 17368 164212
rect 241060 158040 241112 158092
rect 243544 158040 243596 158092
rect 35256 151716 35308 151768
rect 37740 151716 37792 151768
rect 3516 150356 3568 150408
rect 31024 150356 31076 150408
rect 241152 143488 241204 143540
rect 371884 143488 371936 143540
rect 284944 139340 284996 139392
rect 580172 139340 580224 139392
rect 3516 137912 3568 137964
rect 24124 137912 24176 137964
rect 241428 137912 241480 137964
rect 385684 137912 385736 137964
rect 35348 135124 35400 135176
rect 38016 135124 38068 135176
rect 38292 128324 38344 128376
rect 40500 128324 40552 128376
rect 241428 128256 241480 128308
rect 294604 128256 294656 128308
rect 341524 126896 341576 126948
rect 580172 126896 580224 126948
rect 35716 124108 35768 124160
rect 38016 124108 38068 124160
rect 279424 113092 279476 113144
rect 579620 113092 579672 113144
rect 240876 113024 240928 113076
rect 291844 113024 291896 113076
rect 3148 111732 3200 111784
rect 19984 111732 20036 111784
rect 35440 107584 35492 107636
rect 38016 107584 38068 107636
rect 241428 107584 241480 107636
rect 367744 107584 367796 107636
rect 241244 103436 241296 103488
rect 337476 103436 337528 103488
rect 283564 100648 283616 100700
rect 580172 100648 580224 100700
rect 241428 93780 241480 93832
rect 373264 93780 373316 93832
rect 241428 88272 241480 88324
rect 361580 88272 361632 88324
rect 268384 86912 268436 86964
rect 579620 86912 579672 86964
rect 3148 85484 3200 85536
rect 25504 85484 25556 85536
rect 241244 78616 241296 78668
rect 360200 78616 360252 78668
rect 35532 75828 35584 75880
rect 38016 75828 38068 75880
rect 276664 73108 276716 73160
rect 580172 73108 580224 73160
rect 3148 71612 3200 71664
rect 6184 71612 6236 71664
rect 241428 67532 241480 67584
rect 351184 67532 351236 67584
rect 241244 63452 241296 63504
rect 358820 63452 358872 63504
rect 3056 59304 3108 59356
rect 13084 59304 13136 59356
rect 241428 52368 241480 52420
rect 362960 52368 363012 52420
rect 267004 46860 267056 46912
rect 580172 46860 580224 46912
rect 3424 45500 3476 45552
rect 28264 45500 28316 45552
rect 35808 42712 35860 42764
rect 38016 42712 38068 42764
rect 58256 39856 58308 39908
rect 191564 39856 191616 39908
rect 234896 39856 234948 39908
rect 238852 39856 238904 39908
rect 233516 39380 233568 39432
rect 241520 39380 241572 39432
rect 38476 39312 38528 39364
rect 106464 39312 106516 39364
rect 202052 39312 202104 39364
rect 255964 39312 256016 39364
rect 196808 39244 196860 39296
rect 287704 39244 287756 39296
rect 199476 39176 199528 39228
rect 352564 39176 352616 39228
rect 232228 39108 232280 39160
rect 411904 39108 411956 39160
rect 223028 39040 223080 39092
rect 406384 39040 406436 39092
rect 224408 38972 224460 39024
rect 409144 38972 409196 39024
rect 211252 38904 211304 38956
rect 399484 38904 399536 38956
rect 212540 38836 212592 38888
rect 402244 38836 402296 38888
rect 206008 38768 206060 38820
rect 395344 38768 395396 38820
rect 221740 38700 221792 38752
rect 420920 38700 420972 38752
rect 228272 38632 228324 38684
rect 434720 38632 434772 38684
rect 39304 38564 39356 38616
rect 40684 38564 40736 38616
rect 183652 38564 183704 38616
rect 217784 38564 217836 38616
rect 237932 38564 237984 38616
rect 40316 38496 40368 38548
rect 186320 38496 186372 38548
rect 220452 38496 220504 38548
rect 238116 38496 238168 38548
rect 51724 38428 51776 38480
rect 61660 38428 61712 38480
rect 106464 38428 106516 38480
rect 195520 38428 195572 38480
rect 229652 38428 229704 38480
rect 392584 38428 392636 38480
rect 53104 38360 53156 38412
rect 87880 38360 87932 38412
rect 226984 38360 227036 38412
rect 238024 38360 238076 38412
rect 10968 38292 11020 38344
rect 51172 38292 51224 38344
rect 54484 38292 54536 38344
rect 91836 38292 91888 38344
rect 190276 38292 190328 38344
rect 258724 38292 258776 38344
rect 15108 38224 15160 38276
rect 56416 38224 56468 38276
rect 60372 38224 60424 38276
rect 68192 38224 68244 38276
rect 194140 38224 194192 38276
rect 261484 38224 261536 38276
rect 24768 38156 24820 38208
rect 66904 38156 66956 38208
rect 198096 38156 198148 38208
rect 262864 38156 262916 38208
rect 37188 38088 37240 38140
rect 79968 38088 80020 38140
rect 225696 38088 225748 38140
rect 290464 38088 290516 38140
rect 33048 38020 33100 38072
rect 76104 38020 76156 38072
rect 208584 38020 208636 38072
rect 250444 38020 250496 38072
rect 28908 37952 28960 38004
rect 72148 37952 72200 38004
rect 81440 37952 81492 38004
rect 82636 37952 82688 38004
rect 106372 37952 106424 38004
rect 107568 37952 107620 38004
rect 135260 37952 135312 38004
rect 136456 37952 136508 38004
rect 159364 37952 159416 38004
rect 160100 37952 160152 38004
rect 160192 37952 160244 38004
rect 161388 37952 161440 38004
rect 161480 37952 161532 38004
rect 162676 37952 162728 38004
rect 179788 37952 179840 38004
rect 180708 37952 180760 38004
rect 182364 37952 182416 38004
rect 183468 37952 183520 38004
rect 213828 37952 213880 38004
rect 380164 37952 380216 38004
rect 39948 37884 40000 37936
rect 83924 37884 83976 37936
rect 162124 37884 162176 37936
rect 163964 37884 164016 37936
rect 219164 37884 219216 37936
rect 384304 37884 384356 37936
rect 55864 37816 55916 37868
rect 57704 37816 57756 37868
rect 100024 37816 100076 37868
rect 101036 37816 101088 37868
rect 181076 37816 181128 37868
rect 182088 37816 182140 37868
rect 185032 37748 185084 37800
rect 254584 37748 254636 37800
rect 57244 37680 57296 37732
rect 62948 37680 63000 37732
rect 95884 37680 95936 37732
rect 99656 37680 99708 37732
rect 209964 37680 210016 37732
rect 238208 37680 238260 37732
rect 230940 37612 230992 37664
rect 239036 37612 239088 37664
rect 236184 37544 236236 37596
rect 241612 37544 241664 37596
rect 91744 37272 91796 37324
rect 94412 37272 94464 37324
rect 151084 37272 151136 37324
rect 152188 37272 152240 37324
rect 72424 37204 72476 37256
rect 110236 37204 110288 37256
rect 25504 37136 25556 37188
rect 49792 37136 49844 37188
rect 75184 37136 75236 37188
rect 114100 37136 114152 37188
rect 15844 37068 15896 37120
rect 43260 37068 43312 37120
rect 90364 37068 90416 37120
rect 135168 37068 135220 37120
rect 6184 37000 6236 37052
rect 38568 37000 38620 37052
rect 41972 37000 42024 37052
rect 43444 37000 43496 37052
rect 69480 37000 69532 37052
rect 87604 37000 87656 37052
rect 131212 37000 131264 37052
rect 17224 36932 17276 36984
rect 53748 36932 53800 36984
rect 70308 36932 70360 36984
rect 116768 36932 116820 36984
rect 19984 36864 20036 36916
rect 58992 36864 59044 36916
rect 66168 36864 66220 36916
rect 112812 36864 112864 36916
rect 131764 36864 131816 36916
rect 145656 36864 145708 36916
rect 4068 36796 4120 36848
rect 44548 36796 44600 36848
rect 48964 36796 49016 36848
rect 81348 36796 81400 36848
rect 86224 36796 86276 36848
rect 133788 36796 133840 36848
rect 142804 36796 142856 36848
rect 173164 36796 173216 36848
rect 13728 36728 13780 36780
rect 55036 36728 55088 36780
rect 66904 36728 66956 36780
rect 98368 36728 98420 36780
rect 101404 36728 101456 36780
rect 150900 36728 150952 36780
rect 31668 36660 31720 36712
rect 74724 36660 74776 36712
rect 83464 36660 83516 36712
rect 90548 36660 90600 36712
rect 108304 36660 108356 36712
rect 158720 36660 158772 36712
rect 8208 36592 8260 36644
rect 48504 36592 48556 36644
rect 62028 36592 62080 36644
rect 108856 36592 108908 36644
rect 114468 36592 114520 36644
rect 166632 36592 166684 36644
rect 2044 36524 2096 36576
rect 40684 36524 40736 36576
rect 42708 36524 42760 36576
rect 86592 36524 86644 36576
rect 104808 36524 104860 36576
rect 156144 36524 156196 36576
rect 71044 36456 71096 36508
rect 106280 36456 106332 36508
rect 68284 36388 68336 36440
rect 102324 36388 102376 36440
rect 50988 35164 51040 35216
rect 95792 35164 95844 35216
rect 2872 33056 2924 33108
rect 21364 33056 21416 33108
rect 273904 33056 273956 33108
rect 580172 33056 580224 33108
rect 21456 32376 21508 32428
rect 59360 32376 59412 32428
rect 3424 20612 3476 20664
rect 14464 20612 14516 20664
rect 111616 11772 111668 11824
rect 162124 11772 162176 11824
rect 33876 11704 33928 11756
rect 64880 11704 64932 11756
rect 115848 11704 115900 11756
rect 167000 11704 167052 11756
rect 105544 10276 105596 10328
rect 142160 10276 142212 10328
rect 61936 7556 61988 7608
rect 104900 7556 104952 7608
rect 3424 6808 3476 6860
rect 33784 6808 33836 6860
rect 265624 6808 265676 6860
rect 580172 6808 580224 6860
rect 92572 6604 92624 6656
rect 125600 6604 125652 6656
rect 87512 6536 87564 6588
rect 117320 6536 117372 6588
rect 117964 6536 118016 6588
rect 153200 6536 153252 6588
rect 99380 6468 99432 6520
rect 140780 6468 140832 6520
rect 38384 6400 38436 6452
rect 81440 6400 81492 6452
rect 88432 6400 88484 6452
rect 136640 6400 136692 6452
rect 47860 6332 47912 6384
rect 92480 6332 92532 6384
rect 101036 6332 101088 6384
rect 151084 6332 151136 6384
rect 51356 6264 51408 6316
rect 96620 6264 96672 6316
rect 108120 6264 108172 6316
rect 159364 6264 159416 6316
rect 54944 6196 54996 6248
rect 100024 6196 100076 6248
rect 118792 6196 118844 6248
rect 171140 6196 171192 6248
rect 73804 6128 73856 6180
rect 121460 6128 121512 6180
rect 122288 6128 122340 6180
rect 175280 6128 175332 6180
rect 83280 5448 83332 5500
rect 132592 5448 132644 5500
rect 80888 5380 80940 5432
rect 129740 5380 129792 5432
rect 79692 5312 79744 5364
rect 128360 5312 128412 5364
rect 86868 5244 86920 5296
rect 135260 5244 135312 5296
rect 51080 5176 51132 5228
rect 88340 5176 88392 5228
rect 90364 5176 90416 5228
rect 139400 5176 139452 5228
rect 49056 5108 49108 5160
rect 91744 5108 91796 5160
rect 93952 5108 94004 5160
rect 143540 5108 143592 5160
rect 40132 5040 40184 5092
rect 77300 5040 77352 5092
rect 78588 5040 78640 5092
rect 126980 5040 127032 5092
rect 128544 5040 128596 5092
rect 178040 5040 178092 5092
rect 40684 4972 40736 5024
rect 84200 4972 84252 5024
rect 98644 4972 98696 5024
rect 149060 4972 149112 5024
rect 34796 4904 34848 4956
rect 78772 4904 78824 4956
rect 97448 4904 97500 4956
rect 147680 4904 147732 4956
rect 30104 4836 30156 4888
rect 73160 4836 73212 4888
rect 105728 4836 105780 4888
rect 157340 4836 157392 4888
rect 29828 4768 29880 4820
rect 63408 4768 63460 4820
rect 63500 4768 63552 4820
rect 70400 4768 70452 4820
rect 72608 4768 72660 4820
rect 120080 4768 120132 4820
rect 123484 4768 123536 4820
rect 176660 4768 176712 4820
rect 76196 4700 76248 4752
rect 124220 4700 124272 4752
rect 75000 4632 75052 4684
rect 122840 4632 122892 4684
rect 21824 4088 21876 4140
rect 29828 4088 29880 4140
rect 43076 4088 43128 4140
rect 53104 4088 53156 4140
rect 63224 4088 63276 4140
rect 72424 4088 72476 4140
rect 91560 4088 91612 4140
rect 99380 4088 99432 4140
rect 102232 4088 102284 4140
rect 117964 4088 118016 4140
rect 119896 4088 119948 4140
rect 142804 4088 142856 4140
rect 23020 4020 23072 4072
rect 33876 4020 33928 4072
rect 37096 4020 37148 4072
rect 48964 4020 49016 4072
rect 59636 4020 59688 4072
rect 71044 4020 71096 4072
rect 77392 4020 77444 4072
rect 92572 4020 92624 4072
rect 95148 4020 95200 4072
rect 131764 4020 131816 4072
rect 19432 3952 19484 4004
rect 51724 3952 51776 4004
rect 56048 3952 56100 4004
rect 68284 3952 68336 4004
rect 82084 3952 82136 4004
rect 87604 3952 87656 4004
rect 89168 3952 89220 4004
rect 138020 3952 138072 4004
rect 27712 3884 27764 3936
rect 63500 3884 63552 3936
rect 70216 3884 70268 3936
rect 87512 3884 87564 3936
rect 92756 3884 92808 3936
rect 105544 3884 105596 3936
rect 110512 3884 110564 3936
rect 161480 3884 161532 3936
rect 25320 3816 25372 3868
rect 60004 3816 60056 3868
rect 60832 3816 60884 3868
rect 106372 3816 106424 3868
rect 110420 3816 110472 3868
rect 160192 3816 160244 3868
rect 8760 3748 8812 3800
rect 25504 3748 25556 3800
rect 26516 3748 26568 3800
rect 43444 3748 43496 3800
rect 45468 3748 45520 3800
rect 83464 3748 83516 3800
rect 96252 3748 96304 3800
rect 146300 3748 146352 3800
rect 2872 3680 2924 3732
rect 15844 3680 15896 3732
rect 20628 3680 20680 3732
rect 57244 3680 57296 3732
rect 67916 3680 67968 3732
rect 15936 3612 15988 3664
rect 55864 3612 55916 3664
rect 64328 3612 64380 3664
rect 7656 3544 7708 3596
rect 8208 3544 8260 3596
rect 9956 3544 10008 3596
rect 10968 3544 11020 3596
rect 11152 3544 11204 3596
rect 52552 3544 52604 3596
rect 57244 3544 57296 3596
rect 103520 3544 103572 3596
rect 109316 3680 109368 3732
rect 117596 3680 117648 3732
rect 169760 3680 169812 3732
rect 112812 3612 112864 3664
rect 164240 3612 164292 3664
rect 114560 3544 114612 3596
rect 116400 3544 116452 3596
rect 168380 3544 168432 3596
rect 182088 3544 182140 3596
rect 582196 3544 582248 3596
rect 6460 3476 6512 3528
rect 47032 3476 47084 3528
rect 50160 3476 50212 3528
rect 50988 3476 51040 3528
rect 53748 3476 53800 3528
rect 95884 3476 95936 3528
rect 99840 3476 99892 3528
rect 101404 3476 101456 3528
rect 103336 3476 103388 3528
rect 154580 3476 154632 3528
rect 183468 3476 183520 3528
rect 583392 3476 583444 3528
rect 5264 3408 5316 3460
rect 45560 3408 45612 3460
rect 52552 3408 52604 3460
rect 66904 3408 66956 3460
rect 69112 3408 69164 3460
rect 70308 3408 70360 3460
rect 71504 3408 71556 3460
rect 572 3340 624 3392
rect 2044 3340 2096 3392
rect 18236 3340 18288 3392
rect 21456 3340 21508 3392
rect 24216 3340 24268 3392
rect 24768 3340 24820 3392
rect 32404 3340 32456 3392
rect 33048 3340 33100 3392
rect 35992 3340 36044 3392
rect 37188 3340 37240 3392
rect 41880 3340 41932 3392
rect 42708 3340 42760 3392
rect 66720 3340 66772 3392
rect 75184 3340 75236 3392
rect 84476 3340 84528 3392
rect 86224 3340 86276 3392
rect 106924 3408 106976 3460
rect 108304 3408 108356 3460
rect 114008 3408 114060 3460
rect 114468 3408 114520 3460
rect 115204 3408 115256 3460
rect 115848 3408 115900 3460
rect 121092 3408 121144 3460
rect 173900 3408 173952 3460
rect 180708 3408 180760 3460
rect 581000 3408 581052 3460
rect 118884 3340 118936 3392
rect 1676 3272 1728 3324
rect 6184 3272 6236 3324
rect 33600 3272 33652 3324
rect 40132 3272 40184 3324
rect 44272 3272 44324 3324
rect 51080 3272 51132 3324
rect 65524 3272 65576 3324
rect 66168 3272 66220 3324
rect 58440 3136 58492 3188
rect 61936 3136 61988 3188
rect 85672 3136 85724 3188
rect 90272 3136 90324 3188
rect 17040 3068 17092 3120
rect 19984 3068 20036 3120
rect 46664 2932 46716 2984
rect 54484 2932 54536 2984
rect 87972 2932 88024 2984
rect 88432 2932 88484 2984
rect 12348 2864 12400 2916
rect 17224 2864 17276 2916
rect 124680 2796 124732 2848
rect 128544 2796 128596 2848
<< metal2 >>
rect 8086 703520 8198 704960
rect 24278 703520 24390 704960
rect 40470 703520 40582 704960
rect 56754 703520 56866 704960
rect 72946 703520 73058 704960
rect 89138 703520 89250 704960
rect 105422 703520 105534 704960
rect 121614 703520 121726 704960
rect 137806 703520 137918 704960
rect 154090 703520 154202 704960
rect 170282 703520 170394 704960
rect 186474 703520 186586 704960
rect 202758 703520 202870 704960
rect 218072 703582 218836 703610
rect 8128 702434 8156 703520
rect 8128 702406 8248 702434
rect 2778 684312 2834 684321
rect 2778 684247 2834 684256
rect 2792 683670 2820 684247
rect 2780 683664 2832 683670
rect 2780 683606 2832 683612
rect 6184 683664 6236 683670
rect 6184 683606 6236 683612
rect 3422 671256 3478 671265
rect 3422 671191 3478 671200
rect 3330 606112 3386 606121
rect 3330 606047 3386 606056
rect 3344 605878 3372 606047
rect 3332 605872 3384 605878
rect 3332 605814 3384 605820
rect 3330 580000 3386 580009
rect 3330 579935 3386 579944
rect 3344 579698 3372 579935
rect 3332 579692 3384 579698
rect 3332 579634 3384 579640
rect 3330 553888 3386 553897
rect 3330 553823 3386 553832
rect 3344 553450 3372 553823
rect 3332 553444 3384 553450
rect 3332 553386 3384 553392
rect 3330 527912 3386 527921
rect 3330 527847 3386 527856
rect 3344 527202 3372 527847
rect 3332 527196 3384 527202
rect 3332 527138 3384 527144
rect 3330 514856 3386 514865
rect 3330 514791 3332 514800
rect 3384 514791 3386 514800
rect 3332 514762 3384 514768
rect 2870 501800 2926 501809
rect 2870 501735 2926 501744
rect 2884 501022 2912 501735
rect 2872 501016 2924 501022
rect 2872 500958 2924 500964
rect 3330 475688 3386 475697
rect 3330 475623 3386 475632
rect 3344 474774 3372 475623
rect 3332 474768 3384 474774
rect 3332 474710 3384 474716
rect 3330 462632 3386 462641
rect 3330 462567 3386 462576
rect 3344 462398 3372 462567
rect 3332 462392 3384 462398
rect 3332 462334 3384 462340
rect 3330 449576 3386 449585
rect 3330 449511 3386 449520
rect 3344 448594 3372 449511
rect 3332 448588 3384 448594
rect 3332 448530 3384 448536
rect 3146 423600 3202 423609
rect 3146 423535 3202 423544
rect 3160 422346 3188 423535
rect 3148 422340 3200 422346
rect 3148 422282 3200 422288
rect 3332 397520 3384 397526
rect 3330 397488 3332 397497
rect 3384 397488 3386 397497
rect 3330 397423 3386 397432
rect 3330 371376 3386 371385
rect 3330 371311 3386 371320
rect 3344 371278 3372 371311
rect 3332 371272 3384 371278
rect 3332 371214 3384 371220
rect 3054 345400 3110 345409
rect 3054 345335 3110 345344
rect 3068 345098 3096 345335
rect 3056 345092 3108 345098
rect 3056 345034 3108 345040
rect 3436 339386 3464 671191
rect 3514 658200 3570 658209
rect 3514 658135 3570 658144
rect 3528 656946 3556 658135
rect 3516 656940 3568 656946
rect 3516 656882 3568 656888
rect 3516 632120 3568 632126
rect 3514 632088 3516 632097
rect 3568 632088 3570 632097
rect 3514 632023 3570 632032
rect 3514 619168 3570 619177
rect 3514 619103 3570 619112
rect 3424 339380 3476 339386
rect 3424 339322 3476 339328
rect 3528 339318 3556 619103
rect 3606 566944 3662 566953
rect 3606 566879 3662 566888
rect 3516 339312 3568 339318
rect 3516 339254 3568 339260
rect 3620 339182 3648 566879
rect 3698 410544 3754 410553
rect 3698 410479 3754 410488
rect 3608 339176 3660 339182
rect 3608 339118 3660 339124
rect 3422 319288 3478 319297
rect 3422 319223 3478 319232
rect 3436 318850 3464 319223
rect 3424 318844 3476 318850
rect 3424 318786 3476 318792
rect 3422 306232 3478 306241
rect 3422 306167 3478 306176
rect 3436 305046 3464 306167
rect 3424 305040 3476 305046
rect 3424 304982 3476 304988
rect 3422 293176 3478 293185
rect 3422 293111 3478 293120
rect 3436 292602 3464 293111
rect 3424 292596 3476 292602
rect 3424 292538 3476 292544
rect 3054 267200 3110 267209
rect 3054 267135 3110 267144
rect 3068 266422 3096 267135
rect 3056 266416 3108 266422
rect 3056 266358 3108 266364
rect 3422 254144 3478 254153
rect 3422 254079 3478 254088
rect 3436 253978 3464 254079
rect 3424 253972 3476 253978
rect 3424 253914 3476 253920
rect 3712 246430 3740 410479
rect 3790 358456 3846 358465
rect 3790 358391 3846 358400
rect 3804 339114 3832 358391
rect 3792 339108 3844 339114
rect 3792 339050 3844 339056
rect 6196 248130 6224 683606
rect 6184 248124 6236 248130
rect 6184 248066 6236 248072
rect 3700 246424 3752 246430
rect 3700 246366 3752 246372
rect 8220 245138 8248 702406
rect 24320 699718 24348 703520
rect 40512 699718 40540 703520
rect 72988 699718 73016 703520
rect 89180 700330 89208 703520
rect 89168 700324 89220 700330
rect 89168 700266 89220 700272
rect 105464 699718 105492 703520
rect 137848 700398 137876 703520
rect 154132 702434 154160 703520
rect 153212 702406 154160 702434
rect 137836 700392 137888 700398
rect 137836 700334 137888 700340
rect 24308 699712 24360 699718
rect 24308 699654 24360 699660
rect 24768 699712 24820 699718
rect 24768 699654 24820 699660
rect 39856 699712 39908 699718
rect 39856 699654 39908 699660
rect 40500 699712 40552 699718
rect 40500 699654 40552 699660
rect 71780 699712 71832 699718
rect 71780 699654 71832 699660
rect 72976 699712 73028 699718
rect 72976 699654 73028 699660
rect 105452 699712 105504 699718
rect 105452 699654 105504 699660
rect 106188 699712 106240 699718
rect 106188 699654 106240 699660
rect 21364 656940 21416 656946
rect 21364 656882 21416 656888
rect 15844 632120 15896 632126
rect 15844 632062 15896 632068
rect 10324 579692 10376 579698
rect 10324 579634 10376 579640
rect 10336 268462 10364 579634
rect 13084 527196 13136 527202
rect 13084 527138 13136 527144
rect 10324 268456 10376 268462
rect 10324 268398 10376 268404
rect 8208 245132 8260 245138
rect 8208 245074 8260 245080
rect 13096 243846 13124 527138
rect 14464 474768 14516 474774
rect 14464 474710 14516 474716
rect 13084 243840 13136 243846
rect 13084 243782 13136 243788
rect 14476 243710 14504 474710
rect 15856 243914 15884 632062
rect 19984 462392 20036 462398
rect 19984 462334 20036 462340
rect 17224 422340 17276 422346
rect 17224 422282 17276 422288
rect 15844 243908 15896 243914
rect 15844 243850 15896 243856
rect 14464 243704 14516 243710
rect 14464 243646 14516 243652
rect 17236 243642 17264 422282
rect 19996 336190 20024 462334
rect 20076 371272 20128 371278
rect 20076 371214 20128 371220
rect 19984 336184 20036 336190
rect 19984 336126 20036 336132
rect 20088 268394 20116 371214
rect 20076 268388 20128 268394
rect 20076 268330 20128 268336
rect 21376 245614 21404 656882
rect 24780 246838 24808 699654
rect 25504 605872 25556 605878
rect 25504 605814 25556 605820
rect 25516 250918 25544 605814
rect 28264 553444 28316 553450
rect 28264 553386 28316 553392
rect 25504 250912 25556 250918
rect 25504 250854 25556 250860
rect 24768 246832 24820 246838
rect 24768 246774 24820 246780
rect 21364 245608 21416 245614
rect 21364 245550 21416 245556
rect 28276 244866 28304 553386
rect 35164 514820 35216 514826
rect 35164 514762 35216 514768
rect 31024 501016 31076 501022
rect 31024 500958 31076 500964
rect 31036 245546 31064 500958
rect 32404 448588 32456 448594
rect 32404 448530 32456 448536
rect 32416 262954 32444 448530
rect 33784 397520 33836 397526
rect 33784 397462 33836 397468
rect 32404 262948 32456 262954
rect 32404 262890 32456 262896
rect 31024 245540 31076 245546
rect 31024 245482 31076 245488
rect 33796 245478 33824 397462
rect 35176 339454 35204 514762
rect 39764 425740 39816 425746
rect 39764 425682 39816 425688
rect 38382 376952 38438 376961
rect 38382 376887 38438 376896
rect 37554 376000 37610 376009
rect 37554 375935 37610 375944
rect 35624 369912 35676 369918
rect 35624 369854 35676 369860
rect 35256 345092 35308 345098
rect 35256 345034 35308 345040
rect 35164 339448 35216 339454
rect 35164 339390 35216 339396
rect 33784 245472 33836 245478
rect 33784 245414 33836 245420
rect 35268 245274 35296 345034
rect 35348 251864 35400 251870
rect 35348 251806 35400 251812
rect 35256 245268 35308 245274
rect 35256 245210 35308 245216
rect 28264 244860 28316 244866
rect 28264 244802 28316 244808
rect 17224 243636 17276 243642
rect 17224 243578 17276 243584
rect 15936 243500 15988 243506
rect 15936 243442 15988 243448
rect 6184 243160 6236 243166
rect 6184 243102 6236 243108
rect 3424 241664 3476 241670
rect 3424 241606 3476 241612
rect 3436 241097 3464 241606
rect 3422 241088 3478 241097
rect 3422 241023 3478 241032
rect 3424 239216 3476 239222
rect 3424 239158 3476 239164
rect 3332 215280 3384 215286
rect 3332 215222 3384 215228
rect 3344 214985 3372 215222
rect 3330 214976 3386 214985
rect 3330 214911 3386 214920
rect 3056 202836 3108 202842
rect 3056 202778 3108 202784
rect 3068 201929 3096 202778
rect 3054 201920 3110 201929
rect 3054 201855 3110 201864
rect 3240 164212 3292 164218
rect 3240 164154 3292 164160
rect 3252 162897 3280 164154
rect 3238 162888 3294 162897
rect 3238 162823 3294 162832
rect 3148 111784 3200 111790
rect 3148 111726 3200 111732
rect 3160 110673 3188 111726
rect 3146 110664 3202 110673
rect 3146 110599 3202 110608
rect 3436 97617 3464 239158
rect 3516 188896 3568 188902
rect 3514 188864 3516 188873
rect 3568 188864 3570 188873
rect 3514 188799 3570 188808
rect 3516 150408 3568 150414
rect 3516 150350 3568 150356
rect 3528 149841 3556 150350
rect 3514 149832 3570 149841
rect 3514 149767 3570 149776
rect 3516 137964 3568 137970
rect 3516 137906 3568 137912
rect 3528 136785 3556 137906
rect 3514 136776 3570 136785
rect 3514 136711 3570 136720
rect 3422 97608 3478 97617
rect 3422 97543 3478 97552
rect 3148 85536 3200 85542
rect 3148 85478 3200 85484
rect 3160 84697 3188 85478
rect 3146 84688 3202 84697
rect 3146 84623 3202 84632
rect 6196 71670 6224 243102
rect 13084 241596 13136 241602
rect 13084 241538 13136 241544
rect 10324 239352 10376 239358
rect 10324 239294 10376 239300
rect 7564 239284 7616 239290
rect 7564 239226 7616 239232
rect 7576 188902 7604 239226
rect 10336 202842 10364 239294
rect 10324 202836 10376 202842
rect 10324 202778 10376 202784
rect 7564 188896 7616 188902
rect 7564 188838 7616 188844
rect 3148 71664 3200 71670
rect 3146 71632 3148 71641
rect 6184 71664 6236 71670
rect 3200 71632 3202 71641
rect 6184 71606 6236 71612
rect 3146 71567 3202 71576
rect 13096 59362 13124 241538
rect 14464 241528 14516 241534
rect 14464 241470 14516 241476
rect 3056 59356 3108 59362
rect 3056 59298 3108 59304
rect 13084 59356 13136 59362
rect 13084 59298 13136 59304
rect 3068 58585 3096 59298
rect 3054 58576 3110 58585
rect 3054 58511 3110 58520
rect 3424 45552 3476 45558
rect 3422 45520 3424 45529
rect 3476 45520 3478 45529
rect 3422 45455 3478 45464
rect 10968 38344 11020 38350
rect 10968 38286 11020 38292
rect 6184 37052 6236 37058
rect 6184 36994 6236 37000
rect 4068 36848 4120 36854
rect 4068 36790 4120 36796
rect 2044 36576 2096 36582
rect 2044 36518 2096 36524
rect 2056 3398 2084 36518
rect 2872 33108 2924 33114
rect 2872 33050 2924 33056
rect 2884 32473 2912 33050
rect 2870 32464 2926 32473
rect 2870 32399 2926 32408
rect 3424 20664 3476 20670
rect 3424 20606 3476 20612
rect 3436 19417 3464 20606
rect 3422 19408 3478 19417
rect 3422 19343 3478 19352
rect 3424 6860 3476 6866
rect 3424 6802 3476 6808
rect 3436 6497 3464 6802
rect 3422 6488 3478 6497
rect 3422 6423 3478 6432
rect 2872 3732 2924 3738
rect 2872 3674 2924 3680
rect 572 3392 624 3398
rect 572 3334 624 3340
rect 2044 3392 2096 3398
rect 2044 3334 2096 3340
rect 584 480 612 3334
rect 1676 3324 1728 3330
rect 1676 3266 1728 3272
rect 1688 480 1716 3266
rect 2884 480 2912 3674
rect 4080 480 4108 36790
rect 5264 3460 5316 3466
rect 5264 3402 5316 3408
rect 5276 480 5304 3402
rect 6196 3330 6224 36994
rect 8208 36644 8260 36650
rect 8208 36586 8260 36592
rect 8220 3602 8248 36586
rect 8760 3800 8812 3806
rect 8760 3742 8812 3748
rect 7656 3596 7708 3602
rect 7656 3538 7708 3544
rect 8208 3596 8260 3602
rect 8208 3538 8260 3544
rect 6460 3528 6512 3534
rect 6460 3470 6512 3476
rect 6184 3324 6236 3330
rect 6184 3266 6236 3272
rect 6472 480 6500 3470
rect 7668 480 7696 3538
rect 8772 480 8800 3742
rect 10980 3602 11008 38286
rect 13728 36780 13780 36786
rect 13728 36722 13780 36728
rect 13740 6914 13768 36722
rect 14476 20670 14504 241470
rect 15948 215286 15976 243442
rect 28264 243432 28316 243438
rect 28264 243374 28316 243380
rect 17316 243364 17368 243370
rect 17316 243306 17368 243312
rect 15936 215280 15988 215286
rect 15936 215222 15988 215228
rect 17328 164218 17356 243306
rect 19984 243296 20036 243302
rect 19984 243238 20036 243244
rect 17316 164212 17368 164218
rect 17316 164154 17368 164160
rect 19996 111790 20024 243238
rect 21364 243228 21416 243234
rect 21364 243170 21416 243176
rect 19984 111784 20036 111790
rect 19984 111726 20036 111732
rect 15108 38276 15160 38282
rect 15108 38218 15160 38224
rect 14464 20664 14516 20670
rect 14464 20606 14516 20612
rect 15120 6914 15148 38218
rect 15844 37120 15896 37126
rect 15844 37062 15896 37068
rect 13556 6886 13768 6914
rect 14752 6886 15148 6914
rect 9956 3596 10008 3602
rect 9956 3538 10008 3544
rect 10968 3596 11020 3602
rect 10968 3538 11020 3544
rect 11152 3596 11204 3602
rect 11152 3538 11204 3544
rect 9968 480 9996 3538
rect 11164 480 11192 3538
rect 12348 2916 12400 2922
rect 12348 2858 12400 2864
rect 12360 480 12388 2858
rect 13556 480 13584 6886
rect 14752 480 14780 6886
rect 15856 3738 15884 37062
rect 17224 36984 17276 36990
rect 17224 36926 17276 36932
rect 15844 3732 15896 3738
rect 15844 3674 15896 3680
rect 15936 3664 15988 3670
rect 15936 3606 15988 3612
rect 15948 480 15976 3606
rect 17040 3120 17092 3126
rect 17040 3062 17092 3068
rect 17052 480 17080 3062
rect 17236 2922 17264 36926
rect 19984 36916 20036 36922
rect 19984 36858 20036 36864
rect 19432 4004 19484 4010
rect 19432 3946 19484 3952
rect 18236 3392 18288 3398
rect 18236 3334 18288 3340
rect 17224 2916 17276 2922
rect 17224 2858 17276 2864
rect 18248 480 18276 3334
rect 19444 480 19472 3946
rect 19996 3126 20024 36858
rect 21376 33114 21404 243170
rect 25504 239624 25556 239630
rect 25504 239566 25556 239572
rect 24124 239556 24176 239562
rect 24124 239498 24176 239504
rect 24136 137970 24164 239498
rect 24124 137964 24176 137970
rect 24124 137906 24176 137912
rect 25516 85542 25544 239566
rect 25504 85536 25556 85542
rect 25504 85478 25556 85484
rect 28276 45558 28304 243374
rect 35256 242208 35308 242214
rect 35256 242150 35308 242156
rect 33784 239828 33836 239834
rect 33784 239770 33836 239776
rect 31024 239692 31076 239698
rect 31024 239634 31076 239640
rect 31036 150414 31064 239634
rect 31024 150408 31076 150414
rect 31024 150350 31076 150356
rect 28264 45552 28316 45558
rect 28264 45494 28316 45500
rect 24768 38208 24820 38214
rect 24768 38150 24820 38156
rect 21364 33108 21416 33114
rect 21364 33050 21416 33056
rect 21456 32428 21508 32434
rect 21456 32370 21508 32376
rect 20628 3732 20680 3738
rect 20628 3674 20680 3680
rect 19984 3120 20036 3126
rect 19984 3062 20036 3068
rect 20640 480 20668 3674
rect 21468 3398 21496 32370
rect 21824 4140 21876 4146
rect 21824 4082 21876 4088
rect 21456 3392 21508 3398
rect 21456 3334 21508 3340
rect 21836 480 21864 4082
rect 23020 4072 23072 4078
rect 23020 4014 23072 4020
rect 23032 480 23060 4014
rect 24780 3398 24808 38150
rect 33048 38072 33100 38078
rect 33048 38014 33100 38020
rect 28908 38004 28960 38010
rect 28908 37946 28960 37952
rect 25504 37188 25556 37194
rect 25504 37130 25556 37136
rect 25320 3868 25372 3874
rect 25320 3810 25372 3816
rect 24216 3392 24268 3398
rect 24216 3334 24268 3340
rect 24768 3392 24820 3398
rect 24768 3334 24820 3340
rect 24228 480 24256 3334
rect 25332 480 25360 3810
rect 25516 3806 25544 37130
rect 27712 3936 27764 3942
rect 27712 3878 27764 3884
rect 25504 3800 25556 3806
rect 25504 3742 25556 3748
rect 26516 3800 26568 3806
rect 26516 3742 26568 3748
rect 26528 480 26556 3742
rect 27724 480 27752 3878
rect 28920 480 28948 37946
rect 31668 36712 31720 36718
rect 31668 36654 31720 36660
rect 31680 6914 31708 36654
rect 31312 6886 31708 6914
rect 30104 4888 30156 4894
rect 30104 4830 30156 4836
rect 29828 4820 29880 4826
rect 29828 4762 29880 4768
rect 29840 4146 29868 4762
rect 29828 4140 29880 4146
rect 29828 4082 29880 4088
rect 30116 480 30144 4830
rect 31312 480 31340 6886
rect 33060 3398 33088 38014
rect 33796 6866 33824 239770
rect 35268 151774 35296 242150
rect 35256 151768 35308 151774
rect 35256 151710 35308 151716
rect 35360 135182 35388 251806
rect 35532 250708 35584 250714
rect 35532 250650 35584 250656
rect 35440 249076 35492 249082
rect 35440 249018 35492 249024
rect 35348 135176 35400 135182
rect 35348 135118 35400 135124
rect 35452 107642 35480 249018
rect 35440 107636 35492 107642
rect 35440 107578 35492 107584
rect 35544 75886 35572 250650
rect 35636 169522 35664 369854
rect 35808 347880 35860 347886
rect 35808 347822 35860 347828
rect 35716 336116 35768 336122
rect 35716 336058 35768 336064
rect 35624 169516 35676 169522
rect 35624 169458 35676 169464
rect 35728 124166 35756 336058
rect 35716 124160 35768 124166
rect 35716 124102 35768 124108
rect 35532 75880 35584 75886
rect 35532 75822 35584 75828
rect 35820 42770 35848 347822
rect 37096 336320 37148 336326
rect 37096 336262 37148 336268
rect 36636 249688 36688 249694
rect 36636 249630 36688 249636
rect 36544 242276 36596 242282
rect 36544 242218 36596 242224
rect 36556 215801 36584 242218
rect 36542 215792 36598 215801
rect 36542 215727 36598 215736
rect 36648 210497 36676 249630
rect 36820 247580 36872 247586
rect 36820 247522 36872 247528
rect 36728 240848 36780 240854
rect 36728 240790 36780 240796
rect 36634 210488 36690 210497
rect 36634 210423 36690 210432
rect 36740 177993 36768 240790
rect 36832 183433 36860 247522
rect 36912 244792 36964 244798
rect 36912 244734 36964 244740
rect 36818 183424 36874 183433
rect 36818 183359 36874 183368
rect 36726 177984 36782 177993
rect 36726 177919 36782 177928
rect 36924 161673 36952 244734
rect 37004 241052 37056 241058
rect 37004 240994 37056 241000
rect 36910 161664 36966 161673
rect 36910 161599 36966 161608
rect 37016 53417 37044 240994
rect 37108 145489 37136 336262
rect 37188 336252 37240 336258
rect 37188 336194 37240 336200
rect 37094 145480 37150 145489
rect 37094 145415 37150 145424
rect 37200 85921 37228 336194
rect 37568 129169 37596 375935
rect 37922 371104 37978 371113
rect 37922 371039 37978 371048
rect 37936 369918 37964 371039
rect 37924 369912 37976 369918
rect 37924 369854 37976 369860
rect 38198 350024 38254 350033
rect 38198 349959 38254 349968
rect 37646 348120 37702 348129
rect 37646 348055 37702 348064
rect 37660 347886 37688 348055
rect 37648 347880 37700 347886
rect 37648 347822 37700 347828
rect 38212 246498 38240 349959
rect 38396 338978 38424 376887
rect 38750 373824 38806 373833
rect 38750 373759 38806 373768
rect 38474 372872 38530 372881
rect 38474 372807 38530 372816
rect 38384 338972 38436 338978
rect 38384 338914 38436 338920
rect 38384 337068 38436 337074
rect 38384 337010 38436 337016
rect 38200 246492 38252 246498
rect 38200 246434 38252 246440
rect 38108 240984 38160 240990
rect 38108 240926 38160 240932
rect 37740 240916 37792 240922
rect 37740 240858 37792 240864
rect 37752 199617 37780 240858
rect 38016 240032 38068 240038
rect 38016 239974 38068 239980
rect 37924 239964 37976 239970
rect 37924 239906 37976 239912
rect 37832 239896 37884 239902
rect 37832 239838 37884 239844
rect 37738 199608 37794 199617
rect 37738 199543 37794 199552
rect 37844 188737 37872 239838
rect 37830 188728 37886 188737
rect 37830 188663 37886 188672
rect 37832 169516 37884 169522
rect 37832 169458 37884 169464
rect 37740 151768 37792 151774
rect 37740 151710 37792 151716
rect 37752 150929 37780 151710
rect 37738 150920 37794 150929
rect 37738 150855 37794 150864
rect 37554 129160 37610 129169
rect 37554 129095 37610 129104
rect 37844 102105 37872 169458
rect 37936 167113 37964 239906
rect 37922 167104 37978 167113
rect 37922 167039 37978 167048
rect 38028 156369 38056 239974
rect 38014 156360 38070 156369
rect 38014 156295 38070 156304
rect 38016 135176 38068 135182
rect 38016 135118 38068 135124
rect 38028 134609 38056 135118
rect 38014 134600 38070 134609
rect 38014 134535 38070 134544
rect 38016 124160 38068 124166
rect 38016 124102 38068 124108
rect 38028 123865 38056 124102
rect 38014 123856 38070 123865
rect 38014 123791 38070 123800
rect 38120 112985 38148 240926
rect 38292 238196 38344 238202
rect 38292 238138 38344 238144
rect 38200 232824 38252 232830
rect 38200 232766 38252 232772
rect 38106 112976 38162 112985
rect 38106 112911 38162 112920
rect 38016 107636 38068 107642
rect 38016 107578 38068 107584
rect 38028 107545 38056 107578
rect 38014 107536 38070 107545
rect 38014 107471 38070 107480
rect 37830 102096 37886 102105
rect 37830 102031 37886 102040
rect 37186 85912 37242 85921
rect 37186 85847 37242 85856
rect 38016 75880 38068 75886
rect 38016 75822 38068 75828
rect 38028 75041 38056 75822
rect 38014 75032 38070 75041
rect 38014 74967 38070 74976
rect 38212 64297 38240 232766
rect 38304 232014 38332 238138
rect 38292 232008 38344 232014
rect 38292 231950 38344 231956
rect 38292 128376 38344 128382
rect 38292 128318 38344 128324
rect 38304 96801 38332 128318
rect 38290 96792 38346 96801
rect 38290 96727 38346 96736
rect 38396 80481 38424 337010
rect 38382 80472 38438 80481
rect 38382 80407 38438 80416
rect 38198 64288 38254 64297
rect 38198 64223 38254 64232
rect 37002 53408 37058 53417
rect 37002 53343 37058 53352
rect 35808 42764 35860 42770
rect 35808 42706 35860 42712
rect 38016 42764 38068 42770
rect 38016 42706 38068 42712
rect 38028 42673 38056 42706
rect 38014 42664 38070 42673
rect 38014 42599 38070 42608
rect 38488 39370 38516 372807
rect 38658 370016 38714 370025
rect 38658 369951 38714 369960
rect 38566 348392 38622 348401
rect 38566 348327 38622 348336
rect 38580 338094 38608 348327
rect 38568 338088 38620 338094
rect 38568 338030 38620 338036
rect 38580 241466 38608 338030
rect 38672 246362 38700 369951
rect 38764 339046 38792 373759
rect 38842 368248 38898 368257
rect 38842 368183 38898 368192
rect 38752 339040 38804 339046
rect 38752 338982 38804 338988
rect 38752 336048 38804 336054
rect 38752 335990 38804 335996
rect 38660 246356 38712 246362
rect 38660 246298 38712 246304
rect 38568 241460 38620 241466
rect 38568 241402 38620 241408
rect 38660 239148 38712 239154
rect 38660 239090 38712 239096
rect 38568 238740 38620 238746
rect 38568 238682 38620 238688
rect 38580 232121 38608 238682
rect 38566 232112 38622 232121
rect 38566 232047 38622 232056
rect 38568 232008 38620 232014
rect 38568 231950 38620 231956
rect 38580 69737 38608 231950
rect 38566 69728 38622 69737
rect 38566 69663 38622 69672
rect 38672 58857 38700 239090
rect 38764 172553 38792 335990
rect 38856 262886 38884 368183
rect 38844 262880 38896 262886
rect 38844 262822 38896 262828
rect 39580 245064 39632 245070
rect 39580 245006 39632 245012
rect 39304 241460 39356 241466
rect 39304 241402 39356 241408
rect 39396 241460 39448 241466
rect 39396 241402 39448 241408
rect 39120 241392 39172 241398
rect 39120 241334 39172 241340
rect 38844 241120 38896 241126
rect 38844 241062 38896 241068
rect 38750 172544 38806 172553
rect 38750 172479 38806 172488
rect 38856 91361 38884 241062
rect 39028 240168 39080 240174
rect 39028 240110 39080 240116
rect 38936 239420 38988 239426
rect 38936 239362 38988 239368
rect 38948 118425 38976 239362
rect 39040 140049 39068 240110
rect 39132 194177 39160 241334
rect 39212 241324 39264 241330
rect 39212 241266 39264 241272
rect 39224 205057 39252 241266
rect 39210 205048 39266 205057
rect 39210 204983 39266 204992
rect 39118 194168 39174 194177
rect 39118 194103 39174 194112
rect 39026 140040 39082 140049
rect 39026 139975 39082 139984
rect 38934 118416 38990 118425
rect 38934 118351 38990 118360
rect 38842 91352 38898 91361
rect 38842 91287 38898 91296
rect 38658 58848 38714 58857
rect 38658 58783 38714 58792
rect 38566 45520 38622 45529
rect 38566 45455 38622 45464
rect 38476 39364 38528 39370
rect 38476 39306 38528 39312
rect 37188 38140 37240 38146
rect 37188 38082 37240 38088
rect 33876 11756 33928 11762
rect 33876 11698 33928 11704
rect 33784 6860 33836 6866
rect 33784 6802 33836 6808
rect 33888 4078 33916 11698
rect 34796 4956 34848 4962
rect 34796 4898 34848 4904
rect 33876 4072 33928 4078
rect 33876 4014 33928 4020
rect 32404 3392 32456 3398
rect 32404 3334 32456 3340
rect 33048 3392 33100 3398
rect 33048 3334 33100 3340
rect 32416 480 32444 3334
rect 33600 3324 33652 3330
rect 33600 3266 33652 3272
rect 33612 480 33640 3266
rect 34808 480 34836 4898
rect 37096 4072 37148 4078
rect 37096 4014 37148 4020
rect 35992 3392 36044 3398
rect 35992 3334 36044 3340
rect 36004 480 36032 3334
rect 37108 2122 37136 4014
rect 37200 3398 37228 38082
rect 38580 37058 38608 45455
rect 39316 38622 39344 241402
rect 39408 240174 39436 241402
rect 39488 241256 39540 241262
rect 39488 241198 39540 241204
rect 39396 240168 39448 240174
rect 39396 240110 39448 240116
rect 39396 239760 39448 239766
rect 39396 239702 39448 239708
rect 39408 221241 39436 239702
rect 39500 226681 39528 241198
rect 39592 239766 39620 245006
rect 39776 242418 39804 425682
rect 39868 338706 39896 699654
rect 71792 425746 71820 699654
rect 106200 425746 106228 699654
rect 153212 472666 153240 702406
rect 170324 700466 170352 703520
rect 202800 703050 202828 703520
rect 201500 703044 201552 703050
rect 201500 702986 201552 702992
rect 202788 703044 202840 703050
rect 202788 702986 202840 702992
rect 193864 700800 193916 700806
rect 193864 700742 193916 700748
rect 191104 700596 191156 700602
rect 191104 700538 191156 700544
rect 170312 700460 170364 700466
rect 170312 700402 170364 700408
rect 176844 700460 176896 700466
rect 176844 700402 176896 700408
rect 176752 700392 176804 700398
rect 176752 700334 176804 700340
rect 176660 700324 176712 700330
rect 176660 700266 176712 700272
rect 153200 472660 153252 472666
rect 153200 472602 153252 472608
rect 71780 425740 71832 425746
rect 71780 425682 71832 425688
rect 106188 425740 106240 425746
rect 106188 425682 106240 425688
rect 146300 339448 146352 339454
rect 146300 339390 146352 339396
rect 133880 339380 133932 339386
rect 133880 339322 133932 339328
rect 100668 339244 100720 339250
rect 100668 339186 100720 339192
rect 97908 338904 97960 338910
rect 97908 338846 97960 338852
rect 89536 338836 89588 338842
rect 89536 338778 89588 338784
rect 82728 338768 82780 338774
rect 82728 338710 82780 338716
rect 39856 338700 39908 338706
rect 39856 338642 39908 338648
rect 77206 338056 77262 338065
rect 77206 337991 77262 338000
rect 81254 338056 81310 338065
rect 81254 337991 81310 338000
rect 59358 337920 59414 337929
rect 42064 337884 42116 337890
rect 59358 337855 59414 337864
rect 42064 337826 42116 337832
rect 40406 337376 40462 337385
rect 40406 337311 40462 337320
rect 40316 336796 40368 336802
rect 40316 336738 40368 336744
rect 39764 242412 39816 242418
rect 39764 242354 39816 242360
rect 39580 239760 39632 239766
rect 39580 239702 39632 239708
rect 40132 239760 40184 239766
rect 40132 239702 40184 239708
rect 40144 238105 40172 239702
rect 40224 239488 40276 239494
rect 40224 239430 40276 239436
rect 40236 238746 40264 239430
rect 40224 238740 40276 238746
rect 40224 238682 40276 238688
rect 40130 238096 40186 238105
rect 40130 238031 40186 238040
rect 39486 226672 39542 226681
rect 39486 226607 39542 226616
rect 39394 221232 39450 221241
rect 39394 221167 39450 221176
rect 39304 38616 39356 38622
rect 39304 38558 39356 38564
rect 40328 38554 40356 336738
rect 40420 232830 40448 337311
rect 40500 337136 40552 337142
rect 40500 337078 40552 337084
rect 40408 232824 40460 232830
rect 40408 232766 40460 232772
rect 40512 128382 40540 337078
rect 40590 242992 40646 243001
rect 40590 242927 40646 242936
rect 41788 242956 41840 242962
rect 40604 240244 40632 242927
rect 41788 242898 41840 242904
rect 41800 240244 41828 242898
rect 42076 240038 42104 337826
rect 50344 337816 50396 337822
rect 50344 337758 50396 337764
rect 56506 337784 56562 337793
rect 43444 337408 43496 337414
rect 43444 337350 43496 337356
rect 43074 241632 43130 241641
rect 43074 241567 43130 241576
rect 43088 240244 43116 241567
rect 42064 240032 42116 240038
rect 42064 239974 42116 239980
rect 43456 239766 43484 337350
rect 46204 337000 46256 337006
rect 46204 336942 46256 336948
rect 44364 243024 44416 243030
rect 44364 242966 44416 242972
rect 44376 240244 44404 242966
rect 46216 239970 46244 336942
rect 48964 336932 49016 336938
rect 48964 336874 49016 336880
rect 48228 243092 48280 243098
rect 48228 243034 48280 243040
rect 46940 241732 46992 241738
rect 46940 241674 46992 241680
rect 46952 240244 46980 241674
rect 48240 240244 48268 243034
rect 46204 239964 46256 239970
rect 46204 239906 46256 239912
rect 48976 239902 49004 336874
rect 50356 239902 50384 337758
rect 56506 337719 56562 337728
rect 57886 337784 57942 337793
rect 57886 337719 57942 337728
rect 56520 337686 56548 337719
rect 56508 337680 56560 337686
rect 56508 337622 56560 337628
rect 57900 246566 57928 337719
rect 57978 337512 58034 337521
rect 57978 337447 58034 337456
rect 57992 336802 58020 337447
rect 59372 337074 59400 337855
rect 60646 337784 60702 337793
rect 60646 337719 60702 337728
rect 62118 337784 62174 337793
rect 62118 337719 62174 337728
rect 64786 337784 64842 337793
rect 64786 337719 64842 337728
rect 68834 337784 68890 337793
rect 68834 337719 68890 337728
rect 69662 337784 69718 337793
rect 69662 337719 69718 337728
rect 60002 337512 60058 337521
rect 60002 337447 60058 337456
rect 60016 337249 60044 337447
rect 60002 337240 60058 337249
rect 60002 337175 60058 337184
rect 59360 337068 59412 337074
rect 59360 337010 59412 337016
rect 57980 336796 58032 336802
rect 57980 336738 58032 336744
rect 60660 246634 60688 337719
rect 61384 337680 61436 337686
rect 61384 337622 61436 337628
rect 60738 337240 60794 337249
rect 60738 337175 60794 337184
rect 60752 337142 60780 337175
rect 60740 337136 60792 337142
rect 60740 337078 60792 337084
rect 60648 246628 60700 246634
rect 60648 246570 60700 246576
rect 57888 246560 57940 246566
rect 57888 246502 57940 246508
rect 61016 242004 61068 242010
rect 61016 241946 61068 241952
rect 53288 241936 53340 241942
rect 53288 241878 53340 241884
rect 53300 240244 53328 241878
rect 58440 241800 58492 241806
rect 58440 241742 58492 241748
rect 58452 240244 58480 241742
rect 61028 240244 61056 241946
rect 61396 240786 61424 337622
rect 61384 240780 61436 240786
rect 61384 240722 61436 240728
rect 48964 239896 49016 239902
rect 45926 239864 45982 239873
rect 45678 239822 45926 239850
rect 48964 239838 49016 239844
rect 50344 239896 50396 239902
rect 50344 239838 50396 239844
rect 45926 239799 45982 239808
rect 62132 239766 62160 337719
rect 64800 251938 64828 337719
rect 66166 337240 66222 337249
rect 66166 337175 66222 337184
rect 67546 337240 67602 337249
rect 67546 337175 67602 337184
rect 66180 337074 66208 337175
rect 67560 337142 67588 337175
rect 67548 337136 67600 337142
rect 67548 337078 67600 337084
rect 66168 337068 66220 337074
rect 66168 337010 66220 337016
rect 68744 324352 68796 324358
rect 68744 324294 68796 324300
rect 67548 298172 67600 298178
rect 67548 298114 67600 298120
rect 66168 271924 66220 271930
rect 66168 271866 66220 271872
rect 66076 258120 66128 258126
rect 66076 258062 66128 258068
rect 64788 251932 64840 251938
rect 64788 251874 64840 251880
rect 64880 242548 64932 242554
rect 64880 242490 64932 242496
rect 63592 242344 63644 242350
rect 63592 242286 63644 242292
rect 62304 241868 62356 241874
rect 62304 241810 62356 241816
rect 62316 240244 62344 241810
rect 63604 240244 63632 242286
rect 64892 240244 64920 242490
rect 66088 240244 66116 258062
rect 66180 242554 66208 271866
rect 66168 242548 66220 242554
rect 66168 242490 66220 242496
rect 67560 240258 67588 298114
rect 68756 240258 68784 324294
rect 68848 245206 68876 337719
rect 68926 337648 68982 337657
rect 68926 337583 68982 337592
rect 68836 245200 68888 245206
rect 68836 245142 68888 245148
rect 68940 241194 68968 337583
rect 69676 336977 69704 337719
rect 77220 337686 77248 337991
rect 78586 337920 78642 337929
rect 78586 337855 78642 337864
rect 78600 337754 78628 337855
rect 78588 337748 78640 337754
rect 78588 337690 78640 337696
rect 77208 337680 77260 337686
rect 71318 337648 71374 337657
rect 71318 337583 71374 337592
rect 74630 337648 74686 337657
rect 77208 337622 77260 337628
rect 79324 337680 79376 337686
rect 79324 337622 79376 337628
rect 79966 337648 80022 337657
rect 74630 337583 74686 337592
rect 69662 336968 69718 336977
rect 69662 336903 69718 336912
rect 70306 336832 70362 336841
rect 70306 336767 70308 336776
rect 70360 336767 70362 336776
rect 70308 336738 70360 336744
rect 71332 331906 71360 337583
rect 71320 331900 71372 331906
rect 71320 331842 71372 331848
rect 70308 311908 70360 311914
rect 70308 311850 70360 311856
rect 68928 241188 68980 241194
rect 68928 241130 68980 241136
rect 70320 240258 70348 311850
rect 71780 250572 71832 250578
rect 71780 250514 71832 250520
rect 71792 248414 71820 250514
rect 71792 248386 72096 248414
rect 71228 247716 71280 247722
rect 71228 247658 71280 247664
rect 67390 240230 67588 240258
rect 68678 240230 68784 240258
rect 69966 240230 70348 240258
rect 71240 240244 71268 247658
rect 72068 240258 72096 248386
rect 73804 244996 73856 245002
rect 73804 244938 73856 244944
rect 72068 240230 72542 240258
rect 73816 240244 73844 244938
rect 74644 241466 74672 337583
rect 75918 336832 75974 336841
rect 75184 336796 75236 336802
rect 75918 336767 75974 336776
rect 75184 336738 75236 336744
rect 75092 247784 75144 247790
rect 75092 247726 75144 247732
rect 74632 241460 74684 241466
rect 74632 241402 74684 241408
rect 75104 240244 75132 247726
rect 75196 242486 75224 336738
rect 75932 336258 75960 336767
rect 75920 336252 75972 336258
rect 75920 336194 75972 336200
rect 79336 252006 79364 337622
rect 79966 337583 80022 337592
rect 79324 252000 79376 252006
rect 79324 251942 79376 251948
rect 77300 250640 77352 250646
rect 77300 250582 77352 250588
rect 76380 244928 76432 244934
rect 76380 244870 76432 244876
rect 75184 242480 75236 242486
rect 75184 242422 75236 242428
rect 76392 240244 76420 244870
rect 77312 240258 77340 250582
rect 78864 247852 78916 247858
rect 78864 247794 78916 247800
rect 77312 240230 77694 240258
rect 78876 240244 78904 247794
rect 79980 242826 80008 337583
rect 81268 336394 81296 337991
rect 82174 337648 82230 337657
rect 82174 337583 82230 337592
rect 81346 337512 81402 337521
rect 81346 337447 81402 337456
rect 81360 336598 81388 337447
rect 81348 336592 81400 336598
rect 81348 336534 81400 336540
rect 81256 336388 81308 336394
rect 81256 336330 81308 336336
rect 82188 334626 82216 337583
rect 82176 334620 82228 334626
rect 82176 334562 82228 334568
rect 82636 247988 82688 247994
rect 82636 247930 82688 247936
rect 80152 247920 80204 247926
rect 80152 247862 80204 247868
rect 79968 242820 80020 242826
rect 79968 242762 80020 242768
rect 80164 240244 80192 247862
rect 81440 242888 81492 242894
rect 81440 242830 81492 242836
rect 81452 240244 81480 242830
rect 82648 240258 82676 247930
rect 82740 242894 82768 338710
rect 84014 338056 84070 338065
rect 84014 337991 84070 338000
rect 82910 337648 82966 337657
rect 82910 337583 82966 337592
rect 82820 249144 82872 249150
rect 82820 249086 82872 249092
rect 82832 242894 82860 249086
rect 82728 242888 82780 242894
rect 82728 242830 82780 242836
rect 82820 242888 82872 242894
rect 82820 242830 82872 242836
rect 82648 240230 82754 240258
rect 73434 239864 73490 239873
rect 73434 239799 73490 239808
rect 73448 239766 73476 239799
rect 82924 239766 82952 337583
rect 84028 337210 84056 337991
rect 86866 337784 86922 337793
rect 86866 337719 86922 337728
rect 87142 337784 87198 337793
rect 87142 337719 87198 337728
rect 85486 337648 85542 337657
rect 85486 337583 85542 337592
rect 85670 337648 85726 337657
rect 85670 337583 85726 337592
rect 84016 337204 84068 337210
rect 84016 337146 84068 337152
rect 85500 252074 85528 337583
rect 85488 252068 85540 252074
rect 85488 252010 85540 252016
rect 84292 250776 84344 250782
rect 84292 250718 84344 250724
rect 84304 242894 84332 250718
rect 85488 243568 85540 243574
rect 85488 243510 85540 243516
rect 84016 242888 84068 242894
rect 84016 242830 84068 242836
rect 84292 242888 84344 242894
rect 84292 242830 84344 242836
rect 85304 242888 85356 242894
rect 85304 242830 85356 242836
rect 84028 240244 84056 242830
rect 85316 240244 85344 242830
rect 85500 242350 85528 243510
rect 85488 242344 85540 242350
rect 85488 242286 85540 242292
rect 85684 241398 85712 337583
rect 86776 253224 86828 253230
rect 86776 253166 86828 253172
rect 85672 241392 85724 241398
rect 85672 241334 85724 241340
rect 86788 240258 86816 253166
rect 86880 248062 86908 337719
rect 87050 337648 87106 337657
rect 87050 337583 87106 337592
rect 86960 249212 87012 249218
rect 86960 249154 87012 249160
rect 86868 248056 86920 248062
rect 86868 247998 86920 248004
rect 86972 242894 87000 249154
rect 86960 242888 87012 242894
rect 86960 242830 87012 242836
rect 87064 241330 87092 337583
rect 87052 241324 87104 241330
rect 87052 241266 87104 241272
rect 86618 240230 86816 240258
rect 43444 239760 43496 239766
rect 49608 239760 49660 239766
rect 43444 239702 43496 239708
rect 49542 239708 49608 239714
rect 52368 239760 52420 239766
rect 50986 239728 51042 239737
rect 49542 239702 49660 239708
rect 49542 239686 49648 239702
rect 50830 239686 50986 239714
rect 52118 239708 52368 239714
rect 54852 239760 54904 239766
rect 52118 239702 52420 239708
rect 54602 239708 54852 239714
rect 56232 239760 56284 239766
rect 54602 239702 54904 239708
rect 55890 239708 56232 239714
rect 57520 239760 57572 239766
rect 55890 239702 56284 239708
rect 57178 239708 57520 239714
rect 57704 239760 57756 239766
rect 57178 239702 57572 239708
rect 57702 239728 57704 239737
rect 59176 239760 59228 239766
rect 57756 239728 57758 239737
rect 52118 239686 52408 239702
rect 54602 239686 54892 239702
rect 55890 239686 56272 239702
rect 57178 239686 57560 239702
rect 50986 239663 51042 239672
rect 57702 239663 57758 239672
rect 59174 239728 59176 239737
rect 60096 239760 60148 239766
rect 59228 239728 59230 239737
rect 59754 239708 60096 239714
rect 59754 239702 60148 239708
rect 62120 239760 62172 239766
rect 62120 239702 62172 239708
rect 73436 239760 73488 239766
rect 75828 239760 75880 239766
rect 73436 239702 73488 239708
rect 75826 239728 75828 239737
rect 82912 239760 82964 239766
rect 75880 239728 75882 239737
rect 59754 239686 60136 239702
rect 59174 239663 59230 239672
rect 87156 239737 87184 337719
rect 89548 335354 89576 338778
rect 91006 338056 91062 338065
rect 91006 337991 91062 338000
rect 89626 337784 89682 337793
rect 89626 337719 89682 337728
rect 89640 337278 89668 337719
rect 89718 337648 89774 337657
rect 89718 337583 89774 337592
rect 89628 337272 89680 337278
rect 89628 337214 89680 337220
rect 89548 335326 89668 335354
rect 87880 242888 87932 242894
rect 87880 242830 87932 242836
rect 87892 240244 87920 242830
rect 89640 240258 89668 335326
rect 89732 245070 89760 337583
rect 91020 252210 91048 337991
rect 93582 337920 93638 337929
rect 93582 337855 93638 337864
rect 92386 337784 92442 337793
rect 92386 337719 92442 337728
rect 91190 337648 91246 337657
rect 91190 337583 91246 337592
rect 91008 252204 91060 252210
rect 91008 252146 91060 252152
rect 90364 248260 90416 248266
rect 90364 248202 90416 248208
rect 89720 245064 89772 245070
rect 89720 245006 89772 245012
rect 89194 240230 89668 240258
rect 90376 240244 90404 248202
rect 91204 241262 91232 337583
rect 91652 248192 91704 248198
rect 91652 248134 91704 248140
rect 91192 241256 91244 241262
rect 91192 241198 91244 241204
rect 91664 240244 91692 248134
rect 92400 241262 92428 337719
rect 93596 337346 93624 337855
rect 96618 337784 96674 337793
rect 96618 337719 96674 337728
rect 93674 337648 93730 337657
rect 93674 337583 93730 337592
rect 96342 337648 96398 337657
rect 96342 337583 96398 337592
rect 93584 337340 93636 337346
rect 93584 337282 93636 337288
rect 93688 246770 93716 337583
rect 95146 336832 95202 336841
rect 95146 336767 95148 336776
rect 95200 336767 95202 336776
rect 95148 336738 95200 336744
rect 95240 249484 95292 249490
rect 95240 249426 95292 249432
rect 94228 246900 94280 246906
rect 94228 246842 94280 246848
rect 93676 246764 93728 246770
rect 93676 246706 93728 246712
rect 92940 245404 92992 245410
rect 92940 245346 92992 245352
rect 92388 241256 92440 241262
rect 92388 241198 92440 241204
rect 92952 240244 92980 245346
rect 94240 240244 94268 246842
rect 95252 240258 95280 249426
rect 96356 242758 96384 337583
rect 96632 337414 96660 337719
rect 96620 337408 96672 337414
rect 96620 337350 96672 337356
rect 96526 336832 96582 336841
rect 96526 336767 96582 336776
rect 96540 336258 96568 336767
rect 96528 336252 96580 336258
rect 96528 336194 96580 336200
rect 97920 242894 97948 338846
rect 97998 338056 98054 338065
rect 97998 337991 98054 338000
rect 98012 336326 98040 337991
rect 99102 337648 99158 337657
rect 99102 337583 99158 337592
rect 99286 337648 99342 337657
rect 99286 337583 99342 337592
rect 98000 336320 98052 336326
rect 98000 336262 98052 336268
rect 98092 248328 98144 248334
rect 98092 248270 98144 248276
rect 96804 242888 96856 242894
rect 96804 242830 96856 242836
rect 97908 242888 97960 242894
rect 97908 242830 97960 242836
rect 96344 242752 96396 242758
rect 96344 242694 96396 242700
rect 96528 242004 96580 242010
rect 96528 241946 96580 241952
rect 95252 240230 95542 240258
rect 96540 239766 96568 241946
rect 96816 240244 96844 242830
rect 98104 240244 98132 248270
rect 99116 241330 99144 337583
rect 99300 337414 99328 337583
rect 99288 337408 99340 337414
rect 99288 337350 99340 337356
rect 99380 250504 99432 250510
rect 99380 250446 99432 250452
rect 99392 242894 99420 250446
rect 99380 242888 99432 242894
rect 99380 242830 99432 242836
rect 100300 242888 100352 242894
rect 100300 242830 100352 242836
rect 99380 242684 99432 242690
rect 99380 242626 99432 242632
rect 99104 241324 99156 241330
rect 99104 241266 99156 241272
rect 99392 240244 99420 242626
rect 100312 240258 100340 242830
rect 100680 242690 100708 339186
rect 128360 338700 128412 338706
rect 128360 338642 128412 338648
rect 121368 338632 121420 338638
rect 121368 338574 121420 338580
rect 104806 337784 104862 337793
rect 104806 337719 104862 337728
rect 113178 337784 113234 337793
rect 113178 337719 113234 337728
rect 117226 337784 117282 337793
rect 117226 337719 117282 337728
rect 118606 337784 118662 337793
rect 118606 337719 118662 337728
rect 102046 337648 102102 337657
rect 102046 337583 102102 337592
rect 100760 249620 100812 249626
rect 100760 249562 100812 249568
rect 100772 242894 100800 249562
rect 102060 245342 102088 337583
rect 104820 337482 104848 337719
rect 104898 337648 104954 337657
rect 104898 337583 104954 337592
rect 108946 337648 109002 337657
rect 108946 337583 109002 337592
rect 104808 337476 104860 337482
rect 104808 337418 104860 337424
rect 102140 249348 102192 249354
rect 102140 249290 102192 249296
rect 102048 245336 102100 245342
rect 102048 245278 102100 245284
rect 102152 242894 102180 249290
rect 104440 245064 104492 245070
rect 104440 245006 104492 245012
rect 100760 242888 100812 242894
rect 100760 242830 100812 242836
rect 101956 242888 102008 242894
rect 101956 242830 102008 242836
rect 102140 242888 102192 242894
rect 102140 242830 102192 242836
rect 103152 242888 103204 242894
rect 103152 242830 103204 242836
rect 100668 242684 100720 242690
rect 100668 242626 100720 242632
rect 100312 240230 100694 240258
rect 101968 240244 101996 242830
rect 103164 240244 103192 242830
rect 104452 240244 104480 245006
rect 104912 244798 104940 337583
rect 106924 336796 106976 336802
rect 106924 336738 106976 336744
rect 106936 252142 106964 336738
rect 108856 267028 108908 267034
rect 108856 266970 108908 266976
rect 106924 252136 106976 252142
rect 106924 252078 106976 252084
rect 106280 249416 106332 249422
rect 106280 249358 106332 249364
rect 105728 248396 105780 248402
rect 105728 248338 105780 248344
rect 104900 244792 104952 244798
rect 104900 244734 104952 244740
rect 105740 240244 105768 248338
rect 106292 242894 106320 249358
rect 108868 248414 108896 266970
rect 108776 248386 108896 248414
rect 106280 242888 106332 242894
rect 106280 242830 106332 242836
rect 107016 242888 107068 242894
rect 107016 242830 107068 242836
rect 107028 240244 107056 242830
rect 108776 240258 108804 248386
rect 108960 246702 108988 337583
rect 110420 249552 110472 249558
rect 110420 249494 110472 249500
rect 110432 248414 110460 249494
rect 110432 248386 110552 248414
rect 109592 247648 109644 247654
rect 109592 247590 109644 247596
rect 108948 246696 109000 246702
rect 108948 246638 109000 246644
rect 108330 240230 108804 240258
rect 109604 240244 109632 247590
rect 110524 240258 110552 248386
rect 113192 247586 113220 337719
rect 117240 337550 117268 337719
rect 118620 337618 118648 337719
rect 118608 337612 118660 337618
rect 118608 337554 118660 337560
rect 117228 337544 117280 337550
rect 117228 337486 117280 337492
rect 121274 336832 121330 336841
rect 121274 336767 121330 336776
rect 121288 336326 121316 336767
rect 121276 336320 121328 336326
rect 121276 336262 121328 336268
rect 119804 250844 119856 250850
rect 119804 250786 119856 250792
rect 117320 249756 117372 249762
rect 117320 249698 117372 249704
rect 114560 249280 114612 249286
rect 114560 249222 114612 249228
rect 113180 247580 113232 247586
rect 113180 247522 113232 247528
rect 112168 244792 112220 244798
rect 112168 244734 112220 244740
rect 110524 240230 110906 240258
rect 112180 240244 112208 244734
rect 113456 243772 113508 243778
rect 113456 243714 113508 243720
rect 113468 240244 113496 243714
rect 114572 240258 114600 249222
rect 117228 243976 117280 243982
rect 117228 243918 117280 243924
rect 115940 242684 115992 242690
rect 115940 242626 115992 242632
rect 114572 240230 114770 240258
rect 115952 240244 115980 242626
rect 117240 240244 117268 243918
rect 117332 242894 117360 249698
rect 117320 242888 117372 242894
rect 117320 242830 117372 242836
rect 118516 242888 118568 242894
rect 118516 242830 118568 242836
rect 118528 240244 118556 242830
rect 119816 242690 119844 250786
rect 119988 244724 120040 244730
rect 119988 244666 120040 244672
rect 119804 242684 119856 242690
rect 119804 242626 119856 242632
rect 120000 240258 120028 244666
rect 121380 240258 121408 338574
rect 122838 337784 122894 337793
rect 122748 337748 122800 337754
rect 122838 337719 122894 337728
rect 125598 337784 125654 337793
rect 125598 337719 125654 337728
rect 122748 337690 122800 337696
rect 122760 240258 122788 337690
rect 122852 249694 122880 337719
rect 122840 249688 122892 249694
rect 122840 249630 122892 249636
rect 124956 242548 125008 242554
rect 124956 242490 125008 242496
rect 123668 242344 123720 242350
rect 123668 242286 123720 242292
rect 119830 240230 120028 240258
rect 121118 240230 121408 240258
rect 122406 240230 122788 240258
rect 123680 240244 123708 242286
rect 124968 240244 124996 242490
rect 125612 242282 125640 337719
rect 126244 337680 126296 337686
rect 126244 337622 126296 337628
rect 126256 242894 126284 337622
rect 126244 242888 126296 242894
rect 126244 242830 126296 242836
rect 126244 242412 126296 242418
rect 126244 242354 126296 242360
rect 125600 242276 125652 242282
rect 125600 242218 125652 242224
rect 126256 240244 126284 242354
rect 127440 242276 127492 242282
rect 127440 242218 127492 242224
rect 127452 240244 127480 242218
rect 128372 240258 128400 338642
rect 131026 338056 131082 338065
rect 131026 337991 131082 338000
rect 129646 336832 129702 336841
rect 129646 336767 129702 336776
rect 129660 336462 129688 336767
rect 131040 336530 131068 337991
rect 133786 337784 133842 337793
rect 133786 337719 133842 337728
rect 131028 336524 131080 336530
rect 131028 336466 131080 336472
rect 129648 336456 129700 336462
rect 129648 336398 129700 336404
rect 132592 248124 132644 248130
rect 132592 248066 132644 248072
rect 131304 246832 131356 246838
rect 131304 246774 131356 246780
rect 130016 245132 130068 245138
rect 130016 245074 130068 245080
rect 128820 241936 128872 241942
rect 128820 241878 128872 241884
rect 128372 240230 128754 240258
rect 128832 239766 128860 241878
rect 130028 240244 130056 245074
rect 131316 240244 131344 246774
rect 132604 240244 132632 248066
rect 133800 242146 133828 337719
rect 133892 248414 133920 339322
rect 138020 339312 138072 339318
rect 138020 339254 138072 339260
rect 136546 337784 136602 337793
rect 136546 337719 136602 337728
rect 133892 248386 134840 248414
rect 133880 245608 133932 245614
rect 133880 245550 133932 245556
rect 133788 242140 133840 242146
rect 133788 242082 133840 242088
rect 133892 240244 133920 245550
rect 134812 240258 134840 248386
rect 136456 243908 136508 243914
rect 136456 243850 136508 243856
rect 134812 240230 135194 240258
rect 136468 240244 136496 243850
rect 136560 242078 136588 337719
rect 136640 250912 136692 250918
rect 136640 250854 136692 250860
rect 136652 248414 136680 250854
rect 138032 248414 138060 339254
rect 142160 339176 142212 339182
rect 142160 339118 142212 339124
rect 139306 337784 139362 337793
rect 139306 337719 139362 337728
rect 136652 248386 137416 248414
rect 138032 248386 138704 248414
rect 136548 242072 136600 242078
rect 136548 242014 136600 242020
rect 137388 240258 137416 248386
rect 138676 240258 138704 248386
rect 137388 240230 137770 240258
rect 138676 240230 139058 240258
rect 139320 239902 139348 337719
rect 142066 337104 142122 337113
rect 142066 337039 142122 337048
rect 139400 268456 139452 268462
rect 139400 268398 139452 268404
rect 139412 248414 139440 268398
rect 139412 248386 139808 248414
rect 139780 240258 139808 248386
rect 141516 244860 141568 244866
rect 141516 244802 141568 244808
rect 139780 240230 140254 240258
rect 141528 240244 141556 244802
rect 142080 243914 142108 337039
rect 142172 248414 142200 339118
rect 143446 337784 143502 337793
rect 143446 337719 143502 337728
rect 146206 337784 146262 337793
rect 146206 337719 146262 337728
rect 143460 337686 143488 337719
rect 143448 337680 143500 337686
rect 143448 337622 143500 337628
rect 142172 248386 142384 248414
rect 142068 243908 142120 243914
rect 142068 243850 142120 243856
rect 142356 240258 142384 248386
rect 146220 245546 146248 337719
rect 145380 245540 145432 245546
rect 145380 245482 145432 245488
rect 146208 245540 146260 245546
rect 146208 245482 146260 245488
rect 144092 243840 144144 243846
rect 144092 243782 144144 243788
rect 142356 240230 142830 240258
rect 144104 240244 144132 243782
rect 145392 240244 145420 245482
rect 146312 240258 146340 339390
rect 157340 339108 157392 339114
rect 157340 339050 157392 339056
rect 150440 336184 150492 336190
rect 150440 336126 150492 336132
rect 149060 262948 149112 262954
rect 149060 262890 149112 262896
rect 147956 243704 148008 243710
rect 147956 243646 148008 243652
rect 146312 240230 146694 240258
rect 147968 240244 147996 243646
rect 149072 240258 149100 262890
rect 150452 240258 150480 336126
rect 154580 268388 154632 268394
rect 154580 268330 154632 268336
rect 154592 248414 154620 268330
rect 157352 248414 157380 339050
rect 173164 336592 173216 336598
rect 173164 336534 173216 336540
rect 158720 318844 158772 318850
rect 158720 318786 158772 318792
rect 158732 248414 158760 318786
rect 161480 305040 161532 305046
rect 161480 304982 161532 304988
rect 160100 292596 160152 292602
rect 160100 292538 160152 292544
rect 160112 248414 160140 292538
rect 161492 248414 161520 304982
rect 162860 266416 162912 266422
rect 162860 266358 162912 266364
rect 162872 248414 162900 266358
rect 165620 253972 165672 253978
rect 165620 253914 165672 253920
rect 154592 248386 155264 248414
rect 157352 248386 157840 248414
rect 158732 248386 159128 248414
rect 160112 248386 160416 248414
rect 161492 248386 161704 248414
rect 162872 248386 162992 248414
rect 154304 246424 154356 246430
rect 154304 246366 154356 246372
rect 153016 245472 153068 245478
rect 153016 245414 153068 245420
rect 151820 243636 151872 243642
rect 151820 243578 151872 243584
rect 149072 240230 149270 240258
rect 150452 240230 150558 240258
rect 151832 240244 151860 243578
rect 153028 240244 153056 245414
rect 154316 240244 154344 246366
rect 155236 240258 155264 248386
rect 156880 245268 156932 245274
rect 156880 245210 156932 245216
rect 155236 240230 155618 240258
rect 156892 240244 156920 245210
rect 157812 240258 157840 248386
rect 159100 240258 159128 248386
rect 160388 240258 160416 248386
rect 161676 240258 161704 248386
rect 162964 240258 162992 248386
rect 164516 241664 164568 241670
rect 164516 241606 164568 241612
rect 157812 240230 158194 240258
rect 159100 240230 159482 240258
rect 160388 240230 160770 240258
rect 161676 240230 162058 240258
rect 162964 240230 163346 240258
rect 164528 240244 164556 241606
rect 165632 240258 165660 253914
rect 167092 243500 167144 243506
rect 167092 243442 167144 243448
rect 165632 240230 165830 240258
rect 167104 240244 167132 243442
rect 170956 243364 171008 243370
rect 170956 243306 171008 243312
rect 168470 241632 168526 241641
rect 168470 241567 168526 241576
rect 168484 240106 168512 241567
rect 170968 240244 170996 243306
rect 173176 241942 173204 336534
rect 175924 336456 175976 336462
rect 175924 336398 175976 336404
rect 174820 243296 174872 243302
rect 174820 243238 174872 243244
rect 173164 241936 173216 241942
rect 173164 241878 173216 241884
rect 174832 240244 174860 243238
rect 175936 242622 175964 336398
rect 175924 242616 175976 242622
rect 175924 242558 175976 242564
rect 176672 242282 176700 700266
rect 176764 337754 176792 700334
rect 176856 338638 176884 700402
rect 189724 700392 189776 700398
rect 189724 700334 189776 700340
rect 185584 700324 185636 700330
rect 185584 700266 185636 700272
rect 182824 670744 182876 670750
rect 182824 670686 182876 670692
rect 180064 616888 180116 616894
rect 180064 616830 180116 616836
rect 176936 472660 176988 472666
rect 176936 472602 176988 472608
rect 176844 338632 176896 338638
rect 176844 338574 176896 338580
rect 176752 337748 176804 337754
rect 176752 337690 176804 337696
rect 176948 242350 176976 472602
rect 177028 425740 177080 425746
rect 177028 425682 177080 425688
rect 177040 242554 177068 425682
rect 177304 336388 177356 336394
rect 177304 336330 177356 336336
rect 177316 242690 177344 336330
rect 178684 334620 178736 334626
rect 178684 334562 178736 334568
rect 178592 243160 178644 243166
rect 178592 243102 178644 243108
rect 177304 242684 177356 242690
rect 177304 242626 177356 242632
rect 177028 242548 177080 242554
rect 177028 242490 177080 242496
rect 176936 242344 176988 242350
rect 176936 242286 176988 242292
rect 176660 242276 176712 242282
rect 176660 242218 176712 242224
rect 178040 241868 178092 241874
rect 178040 241810 178092 241816
rect 177396 241800 177448 241806
rect 177396 241742 177448 241748
rect 175188 241732 175240 241738
rect 175188 241674 175240 241680
rect 168472 240100 168524 240106
rect 168472 240042 168524 240048
rect 171888 239970 172270 239986
rect 171876 239964 172270 239970
rect 171928 239958 172270 239964
rect 171876 239906 171928 239912
rect 139308 239896 139360 239902
rect 139308 239838 139360 239844
rect 175200 239766 175228 241674
rect 96528 239760 96580 239766
rect 82912 239702 82964 239708
rect 87142 239728 87198 239737
rect 75826 239663 75882 239672
rect 96528 239702 96580 239708
rect 128820 239760 128872 239766
rect 173164 239760 173216 239766
rect 128820 239702 128872 239708
rect 168406 239698 168512 239714
rect 169312 239698 169694 239714
rect 175188 239760 175240 239766
rect 173216 239708 173558 239714
rect 173164 239702 173558 239708
rect 175188 239702 175240 239708
rect 168406 239692 168524 239698
rect 168406 239686 168472 239692
rect 87142 239663 87198 239672
rect 168472 239634 168524 239640
rect 169300 239692 169694 239698
rect 169352 239686 169694 239692
rect 173176 239686 173558 239702
rect 175752 239698 176134 239714
rect 177040 239698 177330 239714
rect 177408 239698 177436 241742
rect 178052 239766 178080 241810
rect 178604 240244 178632 243102
rect 178696 242010 178724 334562
rect 180076 248266 180104 616830
rect 180064 248260 180116 248266
rect 180064 248202 180116 248208
rect 182836 246906 182864 670686
rect 185596 248334 185624 700266
rect 187608 349172 187660 349178
rect 187608 349114 187660 349120
rect 185584 248328 185636 248334
rect 185584 248270 185636 248276
rect 182824 246900 182876 246906
rect 182824 246842 182876 246848
rect 186320 246492 186372 246498
rect 186320 246434 186372 246440
rect 179880 243432 179932 243438
rect 179880 243374 179932 243380
rect 178684 242004 178736 242010
rect 178684 241946 178736 241952
rect 179892 240244 179920 243374
rect 182456 243228 182508 243234
rect 182456 243170 182508 243176
rect 181168 241596 181220 241602
rect 181168 241538 181220 241544
rect 181180 240244 181208 241538
rect 182468 240244 182496 243170
rect 185032 241528 185084 241534
rect 185032 241470 185084 241476
rect 185044 240244 185072 241470
rect 186332 240244 186360 246434
rect 187620 240244 187648 349114
rect 189736 249626 189764 700334
rect 189724 249620 189776 249626
rect 189724 249562 189776 249568
rect 191116 248402 191144 700538
rect 191104 248396 191156 248402
rect 191104 248338 191156 248344
rect 193876 247654 193904 700742
rect 198004 700460 198056 700466
rect 198004 700402 198056 700408
rect 196624 696992 196676 696998
rect 196624 696934 196676 696940
rect 195888 367124 195940 367130
rect 195888 367066 195940 367072
rect 195900 248414 195928 367066
rect 195980 262880 196032 262886
rect 195980 262822 196032 262828
rect 195624 248386 195928 248414
rect 195992 248414 196020 262822
rect 196636 249490 196664 696934
rect 196624 249484 196676 249490
rect 196624 249426 196676 249432
rect 195992 248386 196112 248414
rect 193864 247648 193916 247654
rect 193864 247590 193916 247596
rect 192668 246628 192720 246634
rect 192668 246570 192720 246576
rect 191380 246560 191432 246566
rect 191380 246502 191432 246508
rect 190092 242344 190144 242350
rect 190092 242286 190144 242292
rect 188896 242276 188948 242282
rect 188896 242218 188948 242224
rect 188908 240244 188936 242218
rect 190104 240244 190132 242286
rect 191392 240244 191420 246502
rect 192680 240244 192708 246570
rect 193956 243840 194008 243846
rect 193956 243782 194008 243788
rect 193968 240244 193996 243782
rect 195624 240258 195652 248386
rect 195270 240230 195652 240258
rect 196084 240258 196112 248386
rect 198016 243982 198044 700402
rect 200764 643136 200816 643142
rect 200764 643078 200816 643084
rect 200776 248198 200804 643078
rect 201512 249762 201540 702986
rect 211804 700936 211856 700942
rect 211804 700878 211856 700884
rect 209044 700732 209096 700738
rect 209044 700674 209096 700680
rect 204904 700528 204956 700534
rect 204904 700470 204956 700476
rect 202972 339040 203024 339046
rect 202972 338982 203024 338988
rect 201500 249756 201552 249762
rect 201500 249698 201552 249704
rect 202984 248414 203012 338982
rect 204916 249354 204944 700470
rect 207664 336252 207716 336258
rect 207664 336194 207716 336200
rect 204996 252204 205048 252210
rect 204996 252146 205048 252152
rect 204904 249348 204956 249354
rect 204904 249290 204956 249296
rect 202984 248386 203840 248414
rect 200764 248192 200816 248198
rect 200764 248134 200816 248140
rect 199108 246356 199160 246362
rect 199108 246298 199160 246304
rect 198004 243976 198056 243982
rect 198004 243918 198056 243924
rect 198096 243976 198148 243982
rect 198096 243918 198148 243924
rect 198108 240258 198136 243918
rect 196084 240230 196558 240258
rect 197846 240230 198136 240258
rect 199120 240244 199148 246298
rect 202880 242480 202932 242486
rect 202880 242422 202932 242428
rect 200396 242412 200448 242418
rect 200396 242354 200448 242360
rect 200408 240244 200436 242354
rect 201592 241936 201644 241942
rect 201592 241878 201644 241884
rect 201604 240244 201632 241878
rect 202892 240244 202920 242422
rect 203812 240258 203840 248386
rect 205008 242554 205036 252146
rect 205456 245268 205508 245274
rect 205456 245210 205508 245216
rect 204996 242548 205048 242554
rect 204996 242490 205048 242496
rect 203812 240230 204194 240258
rect 205468 240244 205496 245210
rect 207676 242554 207704 336194
rect 209056 249422 209084 700674
rect 211816 249558 211844 700878
rect 215944 700664 215996 700670
rect 215944 700606 215996 700612
rect 214564 630692 214616 630698
rect 214564 630634 214616 630640
rect 213828 336252 213880 336258
rect 213828 336194 213880 336200
rect 211804 249552 211856 249558
rect 211804 249494 211856 249500
rect 209044 249416 209096 249422
rect 209044 249358 209096 249364
rect 213840 248414 213868 336194
rect 213920 252000 213972 252006
rect 213920 251942 213972 251948
rect 213656 248386 213868 248414
rect 208032 246764 208084 246770
rect 208032 246706 208084 246712
rect 206744 242548 206796 242554
rect 206744 242490 206796 242496
rect 207664 242548 207716 242554
rect 207664 242490 207716 242496
rect 206756 240244 206784 242490
rect 208044 240244 208072 246706
rect 210608 242548 210660 242554
rect 210608 242490 210660 242496
rect 211896 242548 211948 242554
rect 211896 242490 211948 242496
rect 209320 242480 209372 242486
rect 209320 242422 209372 242428
rect 209332 240244 209360 242422
rect 210620 240244 210648 242490
rect 211908 240244 211936 242490
rect 213656 240258 213684 248386
rect 213210 240230 213684 240258
rect 213932 240258 213960 251942
rect 214576 245410 214604 630634
rect 215956 267034 215984 700606
rect 216588 269816 216640 269822
rect 216588 269758 216640 269764
rect 215944 267028 215996 267034
rect 215944 266970 215996 266976
rect 214564 245404 214616 245410
rect 214564 245346 214616 245352
rect 216600 242690 216628 269758
rect 218072 244730 218100 703582
rect 218808 703474 218836 703582
rect 218950 703520 219062 704960
rect 235142 703520 235254 704960
rect 251426 703520 251538 704960
rect 267618 703520 267730 704960
rect 283810 703520 283922 704960
rect 299492 703582 299980 703610
rect 218992 703474 219020 703520
rect 218808 703446 219020 703474
rect 229744 701004 229796 701010
rect 229744 700946 229796 700952
rect 220084 700868 220136 700874
rect 220084 700810 220136 700816
rect 219440 252068 219492 252074
rect 219440 252010 219492 252016
rect 218060 244724 218112 244730
rect 218060 244666 218112 244672
rect 215668 242684 215720 242690
rect 215668 242626 215720 242632
rect 216588 242684 216640 242690
rect 216588 242626 216640 242632
rect 213932 240230 214406 240258
rect 215680 240244 215708 242626
rect 218244 242004 218296 242010
rect 218244 241946 218296 241952
rect 216956 241936 217008 241942
rect 216956 241878 217008 241884
rect 216968 240244 216996 241878
rect 218256 240244 218284 241946
rect 219452 240258 219480 252010
rect 220096 244798 220124 700810
rect 226984 590708 227036 590714
rect 226984 590650 227036 590656
rect 225604 336524 225656 336530
rect 225604 336466 225656 336472
rect 223488 336456 223540 336462
rect 223488 336398 223540 336404
rect 220820 336320 220872 336326
rect 220820 336262 220872 336268
rect 220832 248414 220860 336262
rect 220832 248386 221688 248414
rect 220084 244792 220136 244798
rect 220084 244734 220136 244740
rect 220820 242684 220872 242690
rect 220820 242626 220872 242632
rect 219452 240230 219558 240258
rect 220832 240244 220860 242626
rect 221660 240258 221688 248386
rect 223500 240258 223528 336398
rect 225616 242690 225644 336466
rect 226996 249218 227024 590650
rect 229100 252136 229152 252142
rect 229100 252078 229152 252084
rect 226984 249212 227036 249218
rect 226984 249154 227036 249160
rect 229112 248414 229140 252078
rect 229756 249286 229784 700946
rect 235184 700466 235212 703520
rect 267660 701010 267688 703520
rect 283852 702434 283880 703520
rect 282932 702406 283880 702434
rect 267648 701004 267700 701010
rect 267648 700946 267700 700952
rect 235172 700460 235224 700466
rect 235172 700402 235224 700408
rect 238024 700460 238076 700466
rect 238024 700402 238076 700408
rect 231124 563100 231176 563106
rect 231124 563042 231176 563048
rect 231136 253230 231164 563042
rect 238036 339250 238064 700402
rect 269764 536852 269816 536858
rect 269764 536794 269816 536800
rect 267004 524476 267056 524482
rect 267004 524418 267056 524424
rect 265624 510672 265676 510678
rect 265624 510614 265676 510620
rect 262864 375420 262916 375426
rect 262864 375362 262916 375368
rect 261484 369980 261536 369986
rect 261484 369922 261536 369928
rect 258724 369912 258776 369918
rect 258724 369854 258776 369860
rect 254584 347812 254636 347818
rect 254584 347754 254636 347760
rect 238024 339244 238076 339250
rect 238024 339186 238076 339192
rect 240692 338972 240744 338978
rect 240692 338914 240744 338920
rect 237748 337612 237800 337618
rect 237748 337554 237800 337560
rect 237656 337544 237708 337550
rect 237656 337486 237708 337492
rect 237564 337476 237616 337482
rect 237564 337418 237616 337424
rect 236644 337408 236696 337414
rect 236644 337350 236696 337356
rect 232504 337340 232556 337346
rect 232504 337282 232556 337288
rect 231124 253224 231176 253230
rect 231124 253166 231176 253172
rect 229744 249280 229796 249286
rect 229744 249222 229796 249228
rect 229112 248386 229416 248414
rect 225972 243704 226024 243710
rect 225972 243646 226024 243652
rect 225604 242684 225656 242690
rect 225604 242626 225656 242632
rect 224684 242616 224736 242622
rect 224684 242558 224736 242564
rect 221660 240230 222134 240258
rect 223422 240230 223528 240258
rect 224696 240244 224724 242558
rect 225984 240244 226012 243646
rect 227168 242684 227220 242690
rect 227168 242626 227220 242632
rect 227180 240244 227208 242626
rect 228456 242616 228508 242622
rect 228456 242558 228508 242564
rect 228468 240244 228496 242558
rect 229388 240258 229416 248386
rect 231032 245132 231084 245138
rect 231032 245074 231084 245080
rect 229388 240230 229770 240258
rect 231044 240244 231072 245074
rect 232320 242752 232372 242758
rect 232320 242694 232372 242700
rect 232332 240244 232360 242694
rect 183572 239834 183770 239850
rect 232516 239834 232544 337282
rect 234528 336524 234580 336530
rect 234528 336466 234580 336472
rect 234540 242826 234568 336466
rect 236184 243636 236236 243642
rect 236184 243578 236236 243584
rect 233608 242820 233660 242826
rect 233608 242762 233660 242768
rect 234528 242820 234580 242826
rect 234528 242762 234580 242768
rect 233620 240244 233648 242762
rect 234896 242004 234948 242010
rect 234896 241946 234948 241952
rect 234908 240244 234936 241946
rect 236196 240244 236224 243578
rect 236656 240038 236684 337350
rect 236736 337136 236788 337142
rect 236736 337078 236788 337084
rect 236644 240032 236696 240038
rect 236644 239974 236696 239980
rect 236748 239970 236776 337078
rect 237472 242752 237524 242758
rect 237472 242694 237524 242700
rect 237484 240244 237512 242694
rect 236736 239964 236788 239970
rect 236736 239906 236788 239912
rect 183560 239828 183770 239834
rect 183612 239822 183770 239828
rect 232504 239828 232556 239834
rect 183560 239770 183612 239776
rect 232504 239770 232556 239776
rect 178040 239760 178092 239766
rect 178040 239702 178092 239708
rect 175740 239692 176134 239698
rect 169300 239634 169352 239640
rect 175792 239686 176134 239692
rect 177028 239692 177330 239698
rect 175740 239634 175792 239640
rect 177080 239686 177330 239692
rect 177396 239692 177448 239698
rect 177028 239634 177080 239640
rect 177396 239634 177448 239640
rect 40500 128376 40552 128382
rect 40500 128318 40552 128324
rect 237576 41177 237604 337418
rect 237562 41168 237618 41177
rect 237562 41103 237618 41112
rect 237668 40905 237696 337486
rect 237760 41041 237788 337554
rect 238300 337272 238352 337278
rect 238300 337214 238352 337220
rect 238208 337204 238260 337210
rect 238208 337146 238260 337152
rect 237932 251932 237984 251938
rect 237932 251874 237984 251880
rect 237840 240032 237892 240038
rect 237840 239974 237892 239980
rect 237746 41032 237802 41041
rect 237746 40967 237802 40976
rect 237654 40896 237710 40905
rect 237654 40831 237710 40840
rect 237852 40474 237880 239974
rect 237944 57905 237972 251874
rect 238116 242820 238168 242826
rect 238116 242762 238168 242768
rect 238024 241256 238076 241262
rect 238024 241198 238076 241204
rect 237930 57896 237986 57905
rect 237930 57831 237986 57840
rect 237930 40896 237986 40905
rect 237930 40831 237986 40840
rect 237498 40446 237880 40474
rect 40696 38622 40724 40052
rect 40684 38616 40736 38622
rect 40684 38558 40736 38564
rect 40316 38548 40368 38554
rect 40316 38490 40368 38496
rect 39948 37936 40000 37942
rect 39948 37878 40000 37884
rect 38568 37052 38620 37058
rect 38568 36994 38620 37000
rect 39960 6914 39988 37878
rect 40696 36582 40724 38558
rect 41984 37058 42012 40052
rect 43272 37126 43300 40052
rect 43260 37120 43312 37126
rect 43260 37062 43312 37068
rect 41972 37052 42024 37058
rect 41972 36994 42024 37000
rect 43444 37052 43496 37058
rect 43444 36994 43496 37000
rect 40684 36576 40736 36582
rect 40684 36518 40736 36524
rect 42708 36576 42760 36582
rect 42708 36518 42760 36524
rect 39592 6886 39988 6914
rect 38384 6452 38436 6458
rect 38384 6394 38436 6400
rect 37188 3392 37240 3398
rect 37188 3334 37240 3340
rect 37108 2094 37228 2122
rect 37200 480 37228 2094
rect 38396 480 38424 6394
rect 39592 480 39620 6886
rect 40132 5092 40184 5098
rect 40132 5034 40184 5040
rect 40144 3330 40172 5034
rect 40684 5024 40736 5030
rect 40684 4966 40736 4972
rect 40132 3324 40184 3330
rect 40132 3266 40184 3272
rect 40696 480 40724 4966
rect 42720 3398 42748 36518
rect 43076 4140 43128 4146
rect 43076 4082 43128 4088
rect 41880 3392 41932 3398
rect 41880 3334 41932 3340
rect 42708 3392 42760 3398
rect 42708 3334 42760 3340
rect 41892 480 41920 3334
rect 43088 480 43116 4082
rect 43456 3806 43484 36994
rect 44560 36854 44588 40052
rect 44548 36848 44600 36854
rect 44548 36790 44600 36796
rect 45940 26234 45968 40052
rect 47228 26234 47256 40052
rect 48516 36650 48544 40052
rect 49804 37194 49832 40052
rect 51184 38350 51212 40052
rect 51724 38480 51776 38486
rect 51724 38422 51776 38428
rect 51172 38344 51224 38350
rect 51172 38286 51224 38292
rect 49792 37188 49844 37194
rect 49792 37130 49844 37136
rect 48964 36848 49016 36854
rect 48964 36790 49016 36796
rect 48504 36644 48556 36650
rect 48504 36586 48556 36592
rect 45572 26206 45968 26234
rect 47044 26206 47256 26234
rect 43444 3800 43496 3806
rect 43444 3742 43496 3748
rect 45468 3800 45520 3806
rect 45468 3742 45520 3748
rect 44272 3324 44324 3330
rect 44272 3266 44324 3272
rect 44284 480 44312 3266
rect 45480 480 45508 3742
rect 45572 3466 45600 26206
rect 47044 3534 47072 26206
rect 47860 6384 47912 6390
rect 47860 6326 47912 6332
rect 47032 3528 47084 3534
rect 47032 3470 47084 3476
rect 45560 3460 45612 3466
rect 45560 3402 45612 3408
rect 46664 2984 46716 2990
rect 46664 2926 46716 2932
rect 46676 480 46704 2926
rect 47872 480 47900 6326
rect 48976 4078 49004 36790
rect 50988 35216 51040 35222
rect 50988 35158 51040 35164
rect 49056 5160 49108 5166
rect 49056 5102 49108 5108
rect 48964 4072 49016 4078
rect 48964 4014 49016 4020
rect 49068 2666 49096 5102
rect 51000 3534 51028 35158
rect 51356 6316 51408 6322
rect 51356 6258 51408 6264
rect 51080 5228 51132 5234
rect 51080 5170 51132 5176
rect 50160 3528 50212 3534
rect 50160 3470 50212 3476
rect 50988 3528 51040 3534
rect 50988 3470 51040 3476
rect 48976 2638 49096 2666
rect 48976 480 49004 2638
rect 50172 480 50200 3470
rect 51092 3330 51120 5170
rect 51080 3324 51132 3330
rect 51080 3266 51132 3272
rect 51368 480 51396 6258
rect 51736 4010 51764 38422
rect 52472 35894 52500 40052
rect 53104 38412 53156 38418
rect 53104 38354 53156 38360
rect 52472 35866 52592 35894
rect 51724 4004 51776 4010
rect 51724 3946 51776 3952
rect 52564 3602 52592 35866
rect 53116 4146 53144 38354
rect 53760 36990 53788 40052
rect 54484 38344 54536 38350
rect 54484 38286 54536 38292
rect 53748 36984 53800 36990
rect 53748 36926 53800 36932
rect 53104 4140 53156 4146
rect 53104 4082 53156 4088
rect 52552 3596 52604 3602
rect 52552 3538 52604 3544
rect 53748 3528 53800 3534
rect 53748 3470 53800 3476
rect 52552 3460 52604 3466
rect 52552 3402 52604 3408
rect 52564 480 52592 3402
rect 53760 480 53788 3470
rect 54496 2990 54524 38286
rect 55048 36786 55076 40052
rect 56428 38282 56456 40052
rect 56416 38276 56468 38282
rect 56416 38218 56468 38224
rect 57716 37874 57744 40052
rect 58254 39944 58310 39953
rect 58254 39879 58256 39888
rect 58308 39879 58310 39888
rect 58256 39850 58308 39856
rect 55864 37868 55916 37874
rect 55864 37810 55916 37816
rect 57704 37868 57756 37874
rect 57704 37810 57756 37816
rect 55036 36780 55088 36786
rect 55036 36722 55088 36728
rect 54944 6248 54996 6254
rect 54944 6190 54996 6196
rect 54484 2984 54536 2990
rect 54484 2926 54536 2932
rect 54956 480 54984 6190
rect 55876 3670 55904 37810
rect 57244 37732 57296 37738
rect 57244 37674 57296 37680
rect 56048 4004 56100 4010
rect 56048 3946 56100 3952
rect 55864 3664 55916 3670
rect 55864 3606 55916 3612
rect 56060 480 56088 3946
rect 57256 3738 57284 37674
rect 59004 36922 59032 40052
rect 60292 38026 60320 40052
rect 61672 38486 61700 40052
rect 61660 38480 61712 38486
rect 61660 38422 61712 38428
rect 60372 38276 60424 38282
rect 60372 38218 60424 38224
rect 59372 37998 60320 38026
rect 58992 36916 59044 36922
rect 58992 36858 59044 36864
rect 59372 32434 59400 37998
rect 59360 32428 59412 32434
rect 59360 32370 59412 32376
rect 60384 26234 60412 38218
rect 62960 37738 62988 40052
rect 62948 37732 63000 37738
rect 62948 37674 63000 37680
rect 62028 36644 62080 36650
rect 62028 36586 62080 36592
rect 60016 26206 60412 26234
rect 59636 4072 59688 4078
rect 59636 4014 59688 4020
rect 57244 3732 57296 3738
rect 57244 3674 57296 3680
rect 57244 3596 57296 3602
rect 57244 3538 57296 3544
rect 57256 480 57284 3538
rect 58440 3188 58492 3194
rect 58440 3130 58492 3136
rect 58452 480 58480 3130
rect 59648 480 59676 4014
rect 60016 3874 60044 26206
rect 61936 7608 61988 7614
rect 61936 7550 61988 7556
rect 60004 3868 60056 3874
rect 60004 3810 60056 3816
rect 60832 3868 60884 3874
rect 60832 3810 60884 3816
rect 60844 480 60872 3810
rect 61948 3194 61976 7550
rect 61936 3188 61988 3194
rect 61936 3130 61988 3136
rect 62040 480 62068 36586
rect 64248 26234 64276 40052
rect 65628 26234 65656 40052
rect 66916 38214 66944 40052
rect 68204 38282 68232 40052
rect 68192 38276 68244 38282
rect 68192 38218 68244 38224
rect 66904 38208 66956 38214
rect 66904 38150 66956 38156
rect 69492 37058 69520 40052
rect 69480 37052 69532 37058
rect 69480 36994 69532 37000
rect 70308 36984 70360 36990
rect 70308 36926 70360 36932
rect 66168 36916 66220 36922
rect 66168 36858 66220 36864
rect 63512 26206 64276 26234
rect 64892 26206 65656 26234
rect 63512 4978 63540 26206
rect 64892 11762 64920 26206
rect 64880 11756 64932 11762
rect 64880 11698 64932 11704
rect 63420 4950 63540 4978
rect 63420 4826 63448 4950
rect 63408 4820 63460 4826
rect 63408 4762 63460 4768
rect 63500 4820 63552 4826
rect 63500 4762 63552 4768
rect 63224 4140 63276 4146
rect 63224 4082 63276 4088
rect 63236 480 63264 4082
rect 63512 3942 63540 4762
rect 63500 3936 63552 3942
rect 63500 3878 63552 3884
rect 64328 3664 64380 3670
rect 64328 3606 64380 3612
rect 64340 480 64368 3606
rect 66180 3330 66208 36858
rect 66904 36780 66956 36786
rect 66904 36722 66956 36728
rect 66916 3466 66944 36722
rect 68284 36440 68336 36446
rect 68284 36382 68336 36388
rect 68296 4010 68324 36382
rect 68284 4004 68336 4010
rect 68284 3946 68336 3952
rect 70216 3936 70268 3942
rect 70216 3878 70268 3884
rect 67916 3732 67968 3738
rect 67916 3674 67968 3680
rect 66904 3460 66956 3466
rect 66904 3402 66956 3408
rect 66720 3392 66772 3398
rect 66720 3334 66772 3340
rect 65524 3324 65576 3330
rect 65524 3266 65576 3272
rect 66168 3324 66220 3330
rect 66168 3266 66220 3272
rect 65536 480 65564 3266
rect 66732 480 66760 3334
rect 67928 480 67956 3674
rect 69112 3460 69164 3466
rect 69112 3402 69164 3408
rect 69124 480 69152 3402
rect 70228 1986 70256 3878
rect 70320 3466 70348 36926
rect 70872 26234 70900 40052
rect 72160 38010 72188 40052
rect 72148 38004 72200 38010
rect 72148 37946 72200 37952
rect 72424 37256 72476 37262
rect 72424 37198 72476 37204
rect 71044 36508 71096 36514
rect 71044 36450 71096 36456
rect 70412 26206 70900 26234
rect 70412 4826 70440 26206
rect 70400 4820 70452 4826
rect 70400 4762 70452 4768
rect 71056 4078 71084 36450
rect 72436 4146 72464 37198
rect 73448 26234 73476 40052
rect 74736 36718 74764 40052
rect 76116 38078 76144 40052
rect 76104 38072 76156 38078
rect 76104 38014 76156 38020
rect 75184 37188 75236 37194
rect 75184 37130 75236 37136
rect 74724 36712 74776 36718
rect 74724 36654 74776 36660
rect 73172 26206 73476 26234
rect 73172 4894 73200 26206
rect 73804 6180 73856 6186
rect 73804 6122 73856 6128
rect 73160 4888 73212 4894
rect 73160 4830 73212 4836
rect 72608 4820 72660 4826
rect 72608 4762 72660 4768
rect 72424 4140 72476 4146
rect 72424 4082 72476 4088
rect 71044 4072 71096 4078
rect 71044 4014 71096 4020
rect 70308 3460 70360 3466
rect 70308 3402 70360 3408
rect 71504 3460 71556 3466
rect 71504 3402 71556 3408
rect 70228 1958 70348 1986
rect 70320 480 70348 1958
rect 71516 480 71544 3402
rect 72620 480 72648 4762
rect 73816 480 73844 6122
rect 75000 4684 75052 4690
rect 75000 4626 75052 4632
rect 75012 480 75040 4626
rect 75196 3398 75224 37130
rect 77404 26234 77432 40052
rect 78692 35894 78720 40052
rect 79980 38146 80008 40052
rect 79968 38140 80020 38146
rect 79968 38082 80020 38088
rect 81360 36854 81388 40052
rect 82648 38010 82676 40052
rect 81440 38004 81492 38010
rect 81440 37946 81492 37952
rect 82636 38004 82688 38010
rect 82636 37946 82688 37952
rect 81348 36848 81400 36854
rect 81348 36790 81400 36796
rect 78692 35866 78812 35894
rect 77312 26206 77432 26234
rect 77312 5098 77340 26206
rect 77300 5092 77352 5098
rect 77300 5034 77352 5040
rect 78588 5092 78640 5098
rect 78588 5034 78640 5040
rect 76196 4752 76248 4758
rect 76196 4694 76248 4700
rect 75184 3392 75236 3398
rect 75184 3334 75236 3340
rect 76208 480 76236 4694
rect 77392 4072 77444 4078
rect 77392 4014 77444 4020
rect 77404 480 77432 4014
rect 78600 480 78628 5034
rect 78784 4962 78812 35866
rect 81452 6458 81480 37946
rect 83936 37942 83964 40052
rect 83924 37936 83976 37942
rect 83924 37878 83976 37884
rect 83464 36712 83516 36718
rect 83464 36654 83516 36660
rect 81440 6452 81492 6458
rect 81440 6394 81492 6400
rect 83280 5500 83332 5506
rect 83280 5442 83332 5448
rect 80888 5432 80940 5438
rect 80888 5374 80940 5380
rect 79692 5364 79744 5370
rect 79692 5306 79744 5312
rect 78772 4956 78824 4962
rect 78772 4898 78824 4904
rect 79704 480 79732 5306
rect 80900 480 80928 5374
rect 82084 4004 82136 4010
rect 82084 3946 82136 3952
rect 82096 480 82124 3946
rect 83292 480 83320 5442
rect 83476 3806 83504 36654
rect 85316 26234 85344 40052
rect 86224 36848 86276 36854
rect 86224 36790 86276 36796
rect 84212 26206 85344 26234
rect 84212 5030 84240 26206
rect 84200 5024 84252 5030
rect 84200 4966 84252 4972
rect 83464 3800 83516 3806
rect 83464 3742 83516 3748
rect 86236 3398 86264 36790
rect 86604 36582 86632 40052
rect 87892 38418 87920 40052
rect 87880 38412 87932 38418
rect 87880 38354 87932 38360
rect 87604 37052 87656 37058
rect 87604 36994 87656 37000
rect 86592 36576 86644 36582
rect 86592 36518 86644 36524
rect 87512 6588 87564 6594
rect 87512 6530 87564 6536
rect 86868 5296 86920 5302
rect 86868 5238 86920 5244
rect 84476 3392 84528 3398
rect 84476 3334 84528 3340
rect 86224 3392 86276 3398
rect 86224 3334 86276 3340
rect 84488 480 84516 3334
rect 85672 3188 85724 3194
rect 85672 3130 85724 3136
rect 85684 480 85712 3130
rect 86880 480 86908 5238
rect 87524 3942 87552 6530
rect 87616 4010 87644 36994
rect 89180 26234 89208 40052
rect 90364 37120 90416 37126
rect 90364 37062 90416 37068
rect 88352 26206 89208 26234
rect 88352 5234 88380 26206
rect 90376 6914 90404 37062
rect 90560 36718 90588 40052
rect 91848 38350 91876 40052
rect 91836 38344 91888 38350
rect 91836 38286 91888 38292
rect 91744 37324 91796 37330
rect 91744 37266 91796 37272
rect 90548 36712 90600 36718
rect 90548 36654 90600 36660
rect 90284 6886 90404 6914
rect 88432 6452 88484 6458
rect 88432 6394 88484 6400
rect 88340 5228 88392 5234
rect 88340 5170 88392 5176
rect 87604 4004 87656 4010
rect 87604 3946 87656 3952
rect 87512 3936 87564 3942
rect 87512 3878 87564 3884
rect 88444 2990 88472 6394
rect 89168 4004 89220 4010
rect 89168 3946 89220 3952
rect 87972 2984 88024 2990
rect 87972 2926 88024 2932
rect 88432 2984 88484 2990
rect 88432 2926 88484 2932
rect 87984 480 88012 2926
rect 89180 480 89208 3946
rect 90284 3194 90312 6886
rect 90364 5228 90416 5234
rect 90364 5170 90416 5176
rect 90272 3188 90324 3194
rect 90272 3130 90324 3136
rect 90376 480 90404 5170
rect 91756 5166 91784 37266
rect 93136 26234 93164 40052
rect 94424 37330 94452 40052
rect 94412 37324 94464 37330
rect 94412 37266 94464 37272
rect 95804 35222 95832 40052
rect 95884 37732 95936 37738
rect 95884 37674 95936 37680
rect 95792 35216 95844 35222
rect 95792 35158 95844 35164
rect 92492 26206 93164 26234
rect 92492 6390 92520 26206
rect 92572 6656 92624 6662
rect 92572 6598 92624 6604
rect 92480 6384 92532 6390
rect 92480 6326 92532 6332
rect 91744 5160 91796 5166
rect 91744 5102 91796 5108
rect 91560 4140 91612 4146
rect 91560 4082 91612 4088
rect 91572 480 91600 4082
rect 92584 4078 92612 6598
rect 93952 5160 94004 5166
rect 93952 5102 94004 5108
rect 92572 4072 92624 4078
rect 92572 4014 92624 4020
rect 92756 3936 92808 3942
rect 92756 3878 92808 3884
rect 92768 480 92796 3878
rect 93964 480 93992 5102
rect 95148 4072 95200 4078
rect 95148 4014 95200 4020
rect 95160 480 95188 4014
rect 95896 3534 95924 37674
rect 97092 26234 97120 40052
rect 98380 36786 98408 40052
rect 99668 37738 99696 40052
rect 101048 37874 101076 40052
rect 100024 37868 100076 37874
rect 100024 37810 100076 37816
rect 101036 37868 101088 37874
rect 101036 37810 101088 37816
rect 99656 37732 99708 37738
rect 99656 37674 99708 37680
rect 98368 36780 98420 36786
rect 98368 36722 98420 36728
rect 96632 26206 97120 26234
rect 96632 6322 96660 26206
rect 99380 6520 99432 6526
rect 99380 6462 99432 6468
rect 96620 6316 96672 6322
rect 96620 6258 96672 6264
rect 98644 5024 98696 5030
rect 98644 4966 98696 4972
rect 97448 4956 97500 4962
rect 97448 4898 97500 4904
rect 96252 3800 96304 3806
rect 96252 3742 96304 3748
rect 95884 3528 95936 3534
rect 95884 3470 95936 3476
rect 96264 480 96292 3742
rect 97460 480 97488 4898
rect 98656 480 98684 4966
rect 99392 4146 99420 6462
rect 100036 6254 100064 37810
rect 101404 36780 101456 36786
rect 101404 36722 101456 36728
rect 101036 6384 101088 6390
rect 101036 6326 101088 6332
rect 100024 6248 100076 6254
rect 100024 6190 100076 6196
rect 99380 4140 99432 4146
rect 99380 4082 99432 4088
rect 99840 3528 99892 3534
rect 99840 3470 99892 3476
rect 99852 480 99880 3470
rect 101048 480 101076 6326
rect 101416 3534 101444 36722
rect 102336 36446 102364 40052
rect 102324 36440 102376 36446
rect 102324 36382 102376 36388
rect 103624 26234 103652 40052
rect 104808 36576 104860 36582
rect 104808 36518 104860 36524
rect 103532 26206 103652 26234
rect 102232 4140 102284 4146
rect 102232 4082 102284 4088
rect 101404 3528 101456 3534
rect 101404 3470 101456 3476
rect 102244 480 102272 4082
rect 103532 3602 103560 26206
rect 104820 6914 104848 36518
rect 104912 7614 104940 40052
rect 106292 36514 106320 40052
rect 106464 39364 106516 39370
rect 106464 39306 106516 39312
rect 106476 38486 106504 39306
rect 106464 38480 106516 38486
rect 106464 38422 106516 38428
rect 107580 38010 107608 40052
rect 106372 38004 106424 38010
rect 106372 37946 106424 37952
rect 107568 38004 107620 38010
rect 107568 37946 107620 37952
rect 106280 36508 106332 36514
rect 106280 36450 106332 36456
rect 105544 10328 105596 10334
rect 105544 10270 105596 10276
rect 104900 7608 104952 7614
rect 104900 7550 104952 7556
rect 104544 6886 104848 6914
rect 103520 3596 103572 3602
rect 103520 3538 103572 3544
rect 103336 3528 103388 3534
rect 103336 3470 103388 3476
rect 103348 480 103376 3470
rect 104544 480 104572 6886
rect 105556 3942 105584 10270
rect 105728 4888 105780 4894
rect 105728 4830 105780 4836
rect 105544 3936 105596 3942
rect 105544 3878 105596 3884
rect 105740 480 105768 4830
rect 106384 3874 106412 37946
rect 108304 36712 108356 36718
rect 108304 36654 108356 36660
rect 108120 6316 108172 6322
rect 108120 6258 108172 6264
rect 106372 3868 106424 3874
rect 106372 3810 106424 3816
rect 106924 3460 106976 3466
rect 106924 3402 106976 3408
rect 106936 480 106964 3402
rect 108132 480 108160 6258
rect 108316 3466 108344 36654
rect 108868 36650 108896 40052
rect 110248 37262 110276 40052
rect 110236 37256 110288 37262
rect 110236 37198 110288 37204
rect 108856 36644 108908 36650
rect 108856 36586 108908 36592
rect 111536 26234 111564 40052
rect 112824 36922 112852 40052
rect 114112 37194 114140 40052
rect 114100 37188 114152 37194
rect 114100 37130 114152 37136
rect 112812 36916 112864 36922
rect 112812 36858 112864 36864
rect 114468 36644 114520 36650
rect 114468 36586 114520 36592
rect 110432 26206 111564 26234
rect 110432 3874 110460 26206
rect 111616 11824 111668 11830
rect 111616 11766 111668 11772
rect 110512 3936 110564 3942
rect 110512 3878 110564 3884
rect 110420 3868 110472 3874
rect 110420 3810 110472 3816
rect 109316 3732 109368 3738
rect 109316 3674 109368 3680
rect 108304 3460 108356 3466
rect 108304 3402 108356 3408
rect 109328 480 109356 3674
rect 110524 480 110552 3878
rect 111628 480 111656 11766
rect 112812 3664 112864 3670
rect 112812 3606 112864 3612
rect 112824 480 112852 3606
rect 114480 3466 114508 36586
rect 115492 26234 115520 40052
rect 116780 36990 116808 40052
rect 116768 36984 116820 36990
rect 116768 36926 116820 36932
rect 118068 26234 118096 40052
rect 119356 26234 119384 40052
rect 120736 26234 120764 40052
rect 122024 26234 122052 40052
rect 123312 26234 123340 40052
rect 124600 26234 124628 40052
rect 125980 26234 126008 40052
rect 127268 26234 127296 40052
rect 128556 26234 128584 40052
rect 129936 26234 129964 40052
rect 131224 37058 131252 40052
rect 131212 37052 131264 37058
rect 131212 36994 131264 37000
rect 131764 36916 131816 36922
rect 131764 36858 131816 36864
rect 114572 26206 115520 26234
rect 117332 26206 118096 26234
rect 118896 26206 119384 26234
rect 120092 26206 120764 26234
rect 121472 26206 122052 26234
rect 122852 26206 123340 26234
rect 124232 26206 124628 26234
rect 125612 26206 126008 26234
rect 126992 26206 127296 26234
rect 128372 26206 128584 26234
rect 129752 26206 129964 26234
rect 114572 3602 114600 26206
rect 115848 11756 115900 11762
rect 115848 11698 115900 11704
rect 114560 3596 114612 3602
rect 114560 3538 114612 3544
rect 115860 3466 115888 11698
rect 117332 6594 117360 26206
rect 117320 6588 117372 6594
rect 117320 6530 117372 6536
rect 117964 6588 118016 6594
rect 117964 6530 118016 6536
rect 117976 4146 118004 6530
rect 118792 6248 118844 6254
rect 118792 6190 118844 6196
rect 117964 4140 118016 4146
rect 117964 4082 118016 4088
rect 117596 3732 117648 3738
rect 117596 3674 117648 3680
rect 116400 3596 116452 3602
rect 116400 3538 116452 3544
rect 114008 3460 114060 3466
rect 114008 3402 114060 3408
rect 114468 3460 114520 3466
rect 114468 3402 114520 3408
rect 115204 3460 115256 3466
rect 115204 3402 115256 3408
rect 115848 3460 115900 3466
rect 115848 3402 115900 3408
rect 114020 480 114048 3402
rect 115216 480 115244 3402
rect 116412 480 116440 3538
rect 117608 480 117636 3674
rect 118804 480 118832 6190
rect 118896 3398 118924 26206
rect 120092 4826 120120 26206
rect 121472 6186 121500 26206
rect 121460 6180 121512 6186
rect 121460 6122 121512 6128
rect 122288 6180 122340 6186
rect 122288 6122 122340 6128
rect 120080 4820 120132 4826
rect 120080 4762 120132 4768
rect 119896 4140 119948 4146
rect 119896 4082 119948 4088
rect 118884 3392 118936 3398
rect 118884 3334 118936 3340
rect 119908 480 119936 4082
rect 121092 3460 121144 3466
rect 121092 3402 121144 3408
rect 121104 480 121132 3402
rect 122300 480 122328 6122
rect 122852 4690 122880 26206
rect 123484 4820 123536 4826
rect 123484 4762 123536 4768
rect 122840 4684 122892 4690
rect 122840 4626 122892 4632
rect 123496 480 123524 4762
rect 124232 4758 124260 26206
rect 125612 6662 125640 26206
rect 125600 6656 125652 6662
rect 125600 6598 125652 6604
rect 126992 5098 127020 26206
rect 128372 5370 128400 26206
rect 129752 5438 129780 26206
rect 129740 5432 129792 5438
rect 129740 5374 129792 5380
rect 128360 5364 128412 5370
rect 128360 5306 128412 5312
rect 126980 5092 127032 5098
rect 126980 5034 127032 5040
rect 128544 5092 128596 5098
rect 128544 5034 128596 5040
rect 124220 4752 124272 4758
rect 124220 4694 124272 4700
rect 128556 2854 128584 5034
rect 131776 4078 131804 36858
rect 132512 35894 132540 40052
rect 133800 36854 133828 40052
rect 135180 37126 135208 40052
rect 136468 38010 136496 40052
rect 135260 38004 135312 38010
rect 135260 37946 135312 37952
rect 136456 38004 136508 38010
rect 136456 37946 136508 37952
rect 135168 37120 135220 37126
rect 135168 37062 135220 37068
rect 133788 36848 133840 36854
rect 133788 36790 133840 36796
rect 132512 35866 132632 35894
rect 132604 5506 132632 35866
rect 132592 5500 132644 5506
rect 132592 5442 132644 5448
rect 135272 5302 135300 37946
rect 137756 26234 137784 40052
rect 139044 26234 139072 40052
rect 140424 26234 140452 40052
rect 141712 26234 141740 40052
rect 143000 38026 143028 40052
rect 136652 26206 137784 26234
rect 138032 26206 139072 26234
rect 139412 26206 140452 26234
rect 140792 26206 141740 26234
rect 142172 37998 143028 38026
rect 136652 6458 136680 26206
rect 136640 6452 136692 6458
rect 136640 6394 136692 6400
rect 135260 5296 135312 5302
rect 135260 5238 135312 5244
rect 131764 4072 131816 4078
rect 131764 4014 131816 4020
rect 138032 4010 138060 26206
rect 139412 5234 139440 26206
rect 140792 6526 140820 26206
rect 142172 10334 142200 37998
rect 142804 36848 142856 36854
rect 142804 36790 142856 36796
rect 142160 10328 142212 10334
rect 142160 10270 142212 10276
rect 140780 6520 140832 6526
rect 140780 6462 140832 6468
rect 139400 5228 139452 5234
rect 139400 5170 139452 5176
rect 142816 4146 142844 36790
rect 144288 26234 144316 40052
rect 145668 36922 145696 40052
rect 145656 36916 145708 36922
rect 145656 36858 145708 36864
rect 146956 26234 146984 40052
rect 148244 26234 148272 40052
rect 149532 26234 149560 40052
rect 150912 36786 150940 40052
rect 152200 37330 152228 40052
rect 151084 37324 151136 37330
rect 151084 37266 151136 37272
rect 152188 37324 152240 37330
rect 152188 37266 152240 37272
rect 150900 36780 150952 36786
rect 150900 36722 150952 36728
rect 143552 26206 144316 26234
rect 146312 26206 146984 26234
rect 147692 26206 148272 26234
rect 149072 26206 149560 26234
rect 143552 5166 143580 26206
rect 143540 5160 143592 5166
rect 143540 5102 143592 5108
rect 142804 4140 142856 4146
rect 142804 4082 142856 4088
rect 138020 4004 138072 4010
rect 138020 3946 138072 3952
rect 146312 3806 146340 26206
rect 147692 4962 147720 26206
rect 149072 5030 149100 26206
rect 151096 6390 151124 37266
rect 153488 26234 153516 40052
rect 154868 26234 154896 40052
rect 156156 36582 156184 40052
rect 156144 36576 156196 36582
rect 156144 36518 156196 36524
rect 157444 26234 157472 40052
rect 158732 36718 158760 40052
rect 160112 38010 160140 40052
rect 161400 38010 161428 40052
rect 162688 38010 162716 40052
rect 159364 38004 159416 38010
rect 159364 37946 159416 37952
rect 160100 38004 160152 38010
rect 160100 37946 160152 37952
rect 160192 38004 160244 38010
rect 160192 37946 160244 37952
rect 161388 38004 161440 38010
rect 161388 37946 161440 37952
rect 161480 38004 161532 38010
rect 161480 37946 161532 37952
rect 162676 38004 162728 38010
rect 162676 37946 162728 37952
rect 158720 36712 158772 36718
rect 158720 36654 158772 36660
rect 153212 26206 153516 26234
rect 154592 26206 154896 26234
rect 157352 26206 157472 26234
rect 153212 6594 153240 26206
rect 153200 6588 153252 6594
rect 153200 6530 153252 6536
rect 151084 6384 151136 6390
rect 151084 6326 151136 6332
rect 149060 5024 149112 5030
rect 149060 4966 149112 4972
rect 147680 4956 147732 4962
rect 147680 4898 147732 4904
rect 146300 3800 146352 3806
rect 146300 3742 146352 3748
rect 154592 3534 154620 26206
rect 157352 4894 157380 26206
rect 159376 6322 159404 37946
rect 159364 6316 159416 6322
rect 159364 6258 159416 6264
rect 157340 4888 157392 4894
rect 157340 4830 157392 4836
rect 160204 3874 160232 37946
rect 161492 3942 161520 37946
rect 163976 37942 164004 40052
rect 162124 37936 162176 37942
rect 162124 37878 162176 37884
rect 163964 37936 164016 37942
rect 163964 37878 164016 37884
rect 162136 11830 162164 37878
rect 165356 26234 165384 40052
rect 166644 36650 166672 40052
rect 166632 36644 166684 36650
rect 166632 36586 166684 36592
rect 167932 26234 167960 40052
rect 169220 26234 169248 40052
rect 170600 26234 170628 40052
rect 171888 26234 171916 40052
rect 173176 36854 173204 40052
rect 173164 36848 173216 36854
rect 173164 36790 173216 36796
rect 174556 26234 174584 40052
rect 175844 26234 175872 40052
rect 177132 26234 177160 40052
rect 178420 26234 178448 40052
rect 179800 38010 179828 40052
rect 179788 38004 179840 38010
rect 179788 37946 179840 37952
rect 180708 38004 180760 38010
rect 180708 37946 180760 37952
rect 164252 26206 165384 26234
rect 167012 26206 167960 26234
rect 168392 26206 169248 26234
rect 169772 26206 170628 26234
rect 171152 26206 171916 26234
rect 173912 26206 174584 26234
rect 175292 26206 175872 26234
rect 176672 26206 177160 26234
rect 178052 26206 178448 26234
rect 162124 11824 162176 11830
rect 162124 11766 162176 11772
rect 161480 3936 161532 3942
rect 161480 3878 161532 3884
rect 160192 3868 160244 3874
rect 160192 3810 160244 3816
rect 164252 3670 164280 26206
rect 167012 11762 167040 26206
rect 167000 11756 167052 11762
rect 167000 11698 167052 11704
rect 164240 3664 164292 3670
rect 164240 3606 164292 3612
rect 168392 3602 168420 26206
rect 169772 3738 169800 26206
rect 171152 6254 171180 26206
rect 171140 6248 171192 6254
rect 171140 6190 171192 6196
rect 169760 3732 169812 3738
rect 169760 3674 169812 3680
rect 168380 3596 168432 3602
rect 168380 3538 168432 3544
rect 154580 3528 154632 3534
rect 154580 3470 154632 3476
rect 173912 3466 173940 26206
rect 175292 6186 175320 26206
rect 175280 6180 175332 6186
rect 175280 6122 175332 6128
rect 176672 4826 176700 26206
rect 178052 5098 178080 26206
rect 178040 5092 178092 5098
rect 178040 5034 178092 5040
rect 176660 4820 176712 4826
rect 176660 4762 176712 4768
rect 180720 3466 180748 37946
rect 181088 37874 181116 40052
rect 182376 38010 182404 40052
rect 183664 38622 183692 40052
rect 183652 38616 183704 38622
rect 183652 38558 183704 38564
rect 182364 38004 182416 38010
rect 182364 37946 182416 37952
rect 183468 38004 183520 38010
rect 183468 37946 183520 37952
rect 181076 37868 181128 37874
rect 181076 37810 181128 37816
rect 182088 37868 182140 37874
rect 182088 37810 182140 37816
rect 182100 3602 182128 37810
rect 182088 3596 182140 3602
rect 182088 3538 182140 3544
rect 183480 3534 183508 37946
rect 185044 37806 185072 40052
rect 186332 38554 186360 40052
rect 186320 38548 186372 38554
rect 186320 38490 186372 38496
rect 185032 37800 185084 37806
rect 187620 37777 187648 40052
rect 188908 37913 188936 40052
rect 190288 38350 190316 40052
rect 191576 39914 191604 40052
rect 191564 39908 191616 39914
rect 191564 39850 191616 39856
rect 190276 38344 190328 38350
rect 190276 38286 190328 38292
rect 192864 38049 192892 40052
rect 194152 38282 194180 40052
rect 195532 38486 195560 40052
rect 196820 39302 196848 40052
rect 196808 39296 196860 39302
rect 196808 39238 196860 39244
rect 195520 38480 195572 38486
rect 195520 38422 195572 38428
rect 194140 38276 194192 38282
rect 194140 38218 194192 38224
rect 198108 38214 198136 40052
rect 199488 39234 199516 40052
rect 199476 39228 199528 39234
rect 199476 39170 199528 39176
rect 198096 38208 198148 38214
rect 200776 38185 200804 40052
rect 202064 39370 202092 40052
rect 202052 39364 202104 39370
rect 202052 39306 202104 39312
rect 203352 38593 203380 40052
rect 203338 38584 203394 38593
rect 203338 38519 203394 38528
rect 204732 38321 204760 40052
rect 206020 38826 206048 40052
rect 206008 38820 206060 38826
rect 206008 38762 206060 38768
rect 207308 38457 207336 40052
rect 207294 38448 207350 38457
rect 207294 38383 207350 38392
rect 204718 38312 204774 38321
rect 204718 38247 204774 38256
rect 198096 38150 198148 38156
rect 200762 38176 200818 38185
rect 200762 38111 200818 38120
rect 208596 38078 208624 40052
rect 208584 38072 208636 38078
rect 192850 38040 192906 38049
rect 208584 38014 208636 38020
rect 192850 37975 192906 37984
rect 188894 37904 188950 37913
rect 188894 37839 188950 37848
rect 185032 37742 185084 37748
rect 187606 37768 187662 37777
rect 209976 37738 210004 40052
rect 211264 38962 211292 40052
rect 211252 38956 211304 38962
rect 211252 38898 211304 38904
rect 212552 38894 212580 40052
rect 212540 38888 212592 38894
rect 212540 38830 212592 38836
rect 213840 38010 213868 40052
rect 215220 38593 215248 40052
rect 215206 38584 215262 38593
rect 215206 38519 215262 38528
rect 216508 38457 216536 40052
rect 217796 38622 217824 40052
rect 217784 38616 217836 38622
rect 217784 38558 217836 38564
rect 216494 38448 216550 38457
rect 216494 38383 216550 38392
rect 213828 38004 213880 38010
rect 213828 37946 213880 37952
rect 219176 37942 219204 40052
rect 220464 38554 220492 40052
rect 221752 38758 221780 40052
rect 223040 39098 223068 40052
rect 223028 39092 223080 39098
rect 223028 39034 223080 39040
rect 224420 39030 224448 40052
rect 224408 39024 224460 39030
rect 224408 38966 224460 38972
rect 221740 38752 221792 38758
rect 221740 38694 221792 38700
rect 220452 38548 220504 38554
rect 220452 38490 220504 38496
rect 225708 38146 225736 40052
rect 226996 38418 227024 40052
rect 228284 38690 228312 40052
rect 228272 38684 228324 38690
rect 228272 38626 228324 38632
rect 229664 38486 229692 40052
rect 229652 38480 229704 38486
rect 229652 38422 229704 38428
rect 226984 38412 227036 38418
rect 226984 38354 227036 38360
rect 225696 38140 225748 38146
rect 225696 38082 225748 38088
rect 219164 37936 219216 37942
rect 219164 37878 219216 37884
rect 187606 37703 187662 37712
rect 209964 37732 210016 37738
rect 209964 37674 210016 37680
rect 230952 37670 230980 40052
rect 232240 39166 232268 40052
rect 233528 39438 233556 40052
rect 234908 39914 234936 40052
rect 234896 39908 234948 39914
rect 234896 39850 234948 39856
rect 233516 39432 233568 39438
rect 233516 39374 233568 39380
rect 232228 39160 232280 39166
rect 232228 39102 232280 39108
rect 230940 37664 230992 37670
rect 230940 37606 230992 37612
rect 236196 37602 236224 40052
rect 237944 38622 237972 40831
rect 237932 38616 237984 38622
rect 237932 38558 237984 38564
rect 238036 38418 238064 241198
rect 238128 162353 238156 242762
rect 238220 195974 238248 337146
rect 238312 229090 238340 337214
rect 239404 337068 239456 337074
rect 239404 337010 239456 337016
rect 238760 331900 238812 331906
rect 238760 331842 238812 331848
rect 238300 229084 238352 229090
rect 238300 229026 238352 229032
rect 238208 195968 238260 195974
rect 238208 195910 238260 195916
rect 238114 162344 238170 162353
rect 238114 162279 238170 162288
rect 238772 122641 238800 331842
rect 239312 246696 239364 246702
rect 239312 246638 239364 246644
rect 239220 245336 239272 245342
rect 239220 245278 239272 245284
rect 238944 245200 238996 245206
rect 238944 245142 238996 245148
rect 238852 241324 238904 241330
rect 238852 241266 238904 241272
rect 238758 122632 238814 122641
rect 238758 122567 238814 122576
rect 238206 41168 238262 41177
rect 238206 41103 238262 41112
rect 238114 41032 238170 41041
rect 238114 40967 238170 40976
rect 238128 38554 238156 40967
rect 238116 38548 238168 38554
rect 238116 38490 238168 38496
rect 238024 38412 238076 38418
rect 238024 38354 238076 38360
rect 238220 37738 238248 41103
rect 238864 39914 238892 241266
rect 238956 42537 238984 245142
rect 239128 241188 239180 241194
rect 239128 241130 239180 241136
rect 239036 239896 239088 239902
rect 239036 239838 239088 239844
rect 238942 42528 238998 42537
rect 238942 42463 238998 42472
rect 238852 39908 238904 39914
rect 238852 39850 238904 39856
rect 238208 37732 238260 37738
rect 238208 37674 238260 37680
rect 239048 37670 239076 239838
rect 239140 97617 239168 241130
rect 239232 147665 239260 245278
rect 239324 167657 239352 246638
rect 239416 224806 239444 337010
rect 240600 243908 240652 243914
rect 240600 243850 240652 243856
rect 240508 242888 240560 242894
rect 240508 242830 240560 242836
rect 239496 242140 239548 242146
rect 239496 242082 239548 242088
rect 239404 224800 239456 224806
rect 239404 224742 239456 224748
rect 239508 217705 239536 242082
rect 240140 242072 240192 242078
rect 240140 242014 240192 242020
rect 240152 227769 240180 242014
rect 240416 240780 240468 240786
rect 240416 240722 240468 240728
rect 240324 239964 240376 239970
rect 240324 239906 240376 239912
rect 240138 227760 240194 227769
rect 240138 227695 240194 227704
rect 240232 227044 240284 227050
rect 240232 226986 240284 226992
rect 239494 217696 239550 217705
rect 239494 217631 239550 217640
rect 240140 195968 240192 195974
rect 240140 195910 240192 195916
rect 240152 177721 240180 195910
rect 240138 177712 240194 177721
rect 240138 177647 240194 177656
rect 239310 167648 239366 167657
rect 239310 167583 239366 167592
rect 239218 147656 239274 147665
rect 239218 147591 239274 147600
rect 239126 97608 239182 97617
rect 239126 97543 239182 97552
rect 240244 47433 240272 226986
rect 240336 226098 240364 239906
rect 240428 227050 240456 240722
rect 240416 227044 240468 227050
rect 240416 226986 240468 226992
rect 240324 226092 240376 226098
rect 240324 226034 240376 226040
rect 240324 225888 240376 225894
rect 240324 225830 240376 225836
rect 240336 82521 240364 225830
rect 240416 224800 240468 224806
rect 240416 224742 240468 224748
rect 240322 82512 240378 82521
rect 240322 82447 240378 82456
rect 240428 72457 240456 224742
rect 240520 152697 240548 242830
rect 240612 232801 240640 243850
rect 240598 232792 240654 232801
rect 240598 232727 240654 232736
rect 240600 229084 240652 229090
rect 240600 229026 240652 229032
rect 240612 192681 240640 229026
rect 240598 192672 240654 192681
rect 240598 192607 240654 192616
rect 240506 152688 240562 152697
rect 240506 152623 240562 152632
rect 240704 132569 240732 338914
rect 241520 337680 241572 337686
rect 241520 337622 241572 337628
rect 240876 240032 240928 240038
rect 240876 239974 240928 239980
rect 240888 222737 240916 239974
rect 241152 238740 241204 238746
rect 241152 238682 241204 238688
rect 241164 237833 241192 238682
rect 241150 237824 241206 237833
rect 241150 237759 241206 237768
rect 240874 222728 240930 222737
rect 240874 222663 240930 222672
rect 241244 213920 241296 213926
rect 241244 213862 241296 213868
rect 241256 212809 241284 213862
rect 241242 212800 241298 212809
rect 241242 212735 241298 212744
rect 241428 208344 241480 208350
rect 241428 208286 241480 208292
rect 241440 207777 241468 208286
rect 241426 207768 241482 207777
rect 241426 207703 241482 207712
rect 241428 202836 241480 202842
rect 241428 202778 241480 202784
rect 241440 202745 241468 202778
rect 241426 202736 241482 202745
rect 241426 202671 241482 202680
rect 241428 198688 241480 198694
rect 241428 198630 241480 198636
rect 241440 197713 241468 198630
rect 241426 197704 241482 197713
rect 241426 197639 241482 197648
rect 241428 187672 241480 187678
rect 241426 187640 241428 187649
rect 241480 187640 241482 187649
rect 241426 187575 241482 187584
rect 241428 183524 241480 183530
rect 241428 183466 241480 183472
rect 241440 182753 241468 183466
rect 241426 182744 241482 182753
rect 241426 182679 241482 182688
rect 241244 173664 241296 173670
rect 241244 173606 241296 173612
rect 241256 172689 241284 173606
rect 241242 172680 241298 172689
rect 241242 172615 241298 172624
rect 241060 158092 241112 158098
rect 241060 158034 241112 158040
rect 241072 157593 241100 158034
rect 241058 157584 241114 157593
rect 241058 157519 241114 157528
rect 241152 143540 241204 143546
rect 241152 143482 241204 143488
rect 241164 142633 241192 143482
rect 241150 142624 241206 142633
rect 241150 142559 241206 142568
rect 241428 137964 241480 137970
rect 241428 137906 241480 137912
rect 241440 137601 241468 137906
rect 241426 137592 241482 137601
rect 241426 137527 241482 137536
rect 240690 132560 240746 132569
rect 240690 132495 240746 132504
rect 241428 128308 241480 128314
rect 241428 128250 241480 128256
rect 241440 127673 241468 128250
rect 241426 127664 241482 127673
rect 241426 127599 241482 127608
rect 240876 113076 240928 113082
rect 240876 113018 240928 113024
rect 240888 112577 240916 113018
rect 240874 112568 240930 112577
rect 240874 112503 240930 112512
rect 241428 107636 241480 107642
rect 241428 107578 241480 107584
rect 241440 107545 241468 107578
rect 241426 107536 241482 107545
rect 241426 107471 241482 107480
rect 241244 103488 241296 103494
rect 241244 103430 241296 103436
rect 241256 102513 241284 103430
rect 241242 102504 241298 102513
rect 241242 102439 241298 102448
rect 241428 93832 241480 93838
rect 241428 93774 241480 93780
rect 241440 92585 241468 93774
rect 241426 92576 241482 92585
rect 241426 92511 241482 92520
rect 241428 88324 241480 88330
rect 241428 88266 241480 88272
rect 241440 87553 241468 88266
rect 241426 87544 241482 87553
rect 241426 87479 241482 87488
rect 241244 78668 241296 78674
rect 241244 78610 241296 78616
rect 241256 77489 241284 78610
rect 241242 77480 241298 77489
rect 241242 77415 241298 77424
rect 240414 72448 240470 72457
rect 240414 72383 240470 72392
rect 241428 67584 241480 67590
rect 241426 67552 241428 67561
rect 241480 67552 241482 67561
rect 241426 67487 241482 67496
rect 241244 63504 241296 63510
rect 241244 63446 241296 63452
rect 241256 62529 241284 63446
rect 241242 62520 241298 62529
rect 241242 62455 241298 62464
rect 241426 52456 241482 52465
rect 241426 52391 241428 52400
rect 241480 52391 241482 52400
rect 241428 52362 241480 52368
rect 240230 47424 240286 47433
rect 240230 47359 240286 47368
rect 241532 39438 241560 337622
rect 249064 337136 249116 337142
rect 249064 337078 249116 337084
rect 243544 336388 243596 336394
rect 243544 336330 243596 336336
rect 241704 248056 241756 248062
rect 241704 247998 241756 248004
rect 241612 245540 241664 245546
rect 241612 245482 241664 245488
rect 241520 39432 241572 39438
rect 241520 39374 241572 39380
rect 239036 37664 239088 37670
rect 239036 37606 239088 37612
rect 241624 37602 241652 245482
rect 241716 117609 241744 247998
rect 243556 158098 243584 336330
rect 244924 336320 244976 336326
rect 244924 336262 244976 336268
rect 244936 173670 244964 336262
rect 247684 336184 247736 336190
rect 247684 336126 247736 336132
rect 247696 242010 247724 336126
rect 249076 243982 249104 337078
rect 251824 337068 251876 337074
rect 251824 337010 251876 337016
rect 250444 336592 250496 336598
rect 250444 336534 250496 336540
rect 249064 243976 249116 243982
rect 249064 243918 249116 243924
rect 247684 242004 247736 242010
rect 247684 241946 247736 241952
rect 244924 173664 244976 173670
rect 244924 173606 244976 173612
rect 243544 158092 243596 158098
rect 243544 158034 243596 158040
rect 241702 117600 241758 117609
rect 241702 117535 241758 117544
rect 250456 38078 250484 336534
rect 251836 213926 251864 337010
rect 251824 213920 251876 213926
rect 251824 213862 251876 213868
rect 250444 38072 250496 38078
rect 250444 38014 250496 38020
rect 254596 37806 254624 347754
rect 255964 337204 256016 337210
rect 255964 337146 256016 337152
rect 255976 39370 256004 337146
rect 255964 39364 256016 39370
rect 255964 39306 256016 39312
rect 258736 38350 258764 369854
rect 258724 38344 258776 38350
rect 258724 38286 258776 38292
rect 261496 38282 261524 369922
rect 261484 38276 261536 38282
rect 261484 38218 261536 38224
rect 262876 38214 262904 375362
rect 265636 247994 265664 510614
rect 267016 250782 267044 524418
rect 268384 484424 268436 484430
rect 268384 484366 268436 484372
rect 267004 250776 267056 250782
rect 267004 250718 267056 250724
rect 265624 247988 265676 247994
rect 265624 247930 265676 247936
rect 268396 247926 268424 484366
rect 269776 249150 269804 536794
rect 282932 250850 282960 702406
rect 294604 376780 294656 376786
rect 294604 376722 294656 376728
rect 291844 372632 291896 372638
rect 291844 372574 291896 372580
rect 287704 337272 287756 337278
rect 287704 337214 287756 337220
rect 282920 250844 282972 250850
rect 282920 250786 282972 250792
rect 269764 249144 269816 249150
rect 269764 249086 269816 249092
rect 268384 247920 268436 247926
rect 268384 247862 268436 247868
rect 268384 243092 268436 243098
rect 268384 243034 268436 243040
rect 267004 243024 267056 243030
rect 265622 242992 265678 243001
rect 267004 242966 267056 242972
rect 265622 242927 265678 242936
rect 262864 38208 262916 38214
rect 262864 38150 262916 38156
rect 254584 37800 254636 37806
rect 254584 37742 254636 37748
rect 236184 37596 236236 37602
rect 236184 37538 236236 37544
rect 241612 37596 241664 37602
rect 241612 37538 241664 37544
rect 265636 6866 265664 242927
rect 267016 46918 267044 242966
rect 268396 86970 268424 243034
rect 273904 242956 273956 242962
rect 273904 242898 273956 242904
rect 272524 239148 272576 239154
rect 272524 239090 272576 239096
rect 269764 239080 269816 239086
rect 269764 239022 269816 239028
rect 269776 167006 269804 239022
rect 272536 206990 272564 239090
rect 272524 206984 272576 206990
rect 272524 206926 272576 206932
rect 269764 167000 269816 167006
rect 269764 166942 269816 166948
rect 268384 86964 268436 86970
rect 268384 86906 268436 86912
rect 267004 46912 267056 46918
rect 267004 46854 267056 46860
rect 273916 33114 273944 242898
rect 280804 239012 280856 239018
rect 280804 238954 280856 238960
rect 279424 238944 279476 238950
rect 276662 238912 276718 238921
rect 279424 238886 279476 238892
rect 276662 238847 276718 238856
rect 276676 73166 276704 238847
rect 279436 113150 279464 238886
rect 280816 193186 280844 238954
rect 284944 238876 284996 238882
rect 284944 238818 284996 238824
rect 283562 238776 283618 238785
rect 283562 238711 283618 238720
rect 280804 193180 280856 193186
rect 280804 193122 280856 193128
rect 279424 113144 279476 113150
rect 279424 113086 279476 113092
rect 283576 100706 283604 238711
rect 284956 139398 284984 238818
rect 285680 204944 285732 204950
rect 285680 204886 285732 204892
rect 285692 202842 285720 204886
rect 285680 202836 285732 202842
rect 285680 202778 285732 202784
rect 285680 185632 285732 185638
rect 285680 185574 285732 185580
rect 285692 183530 285720 185574
rect 285680 183524 285732 183530
rect 285680 183466 285732 183472
rect 284944 139392 284996 139398
rect 284944 139334 284996 139340
rect 283564 100700 283616 100706
rect 283564 100642 283616 100648
rect 276664 73160 276716 73166
rect 276664 73102 276716 73108
rect 287716 39302 287744 337214
rect 290464 336660 290516 336666
rect 290464 336602 290516 336608
rect 287704 39296 287756 39302
rect 287704 39238 287756 39244
rect 290476 38146 290504 336602
rect 291856 113082 291884 372574
rect 294616 128314 294644 376722
rect 299492 243778 299520 703582
rect 299952 703474 299980 703582
rect 300094 703520 300206 704960
rect 316286 703520 316398 704960
rect 332478 703520 332590 704960
rect 348762 703520 348874 704960
rect 364954 703520 365066 704960
rect 381146 703520 381258 704960
rect 397430 703520 397542 704960
rect 413622 703520 413734 704960
rect 429814 703520 429926 704960
rect 446098 703520 446210 704960
rect 462290 703520 462402 704960
rect 478482 703520 478594 704960
rect 494766 703520 494878 704960
rect 510958 703520 511070 704960
rect 527150 703520 527262 704960
rect 543434 703520 543546 704960
rect 559626 703520 559738 704960
rect 575818 703520 575930 704960
rect 300136 703474 300164 703520
rect 299952 703446 300164 703474
rect 332520 700942 332548 703520
rect 332508 700936 332560 700942
rect 332508 700878 332560 700884
rect 348804 700874 348832 703520
rect 348792 700868 348844 700874
rect 348792 700810 348844 700816
rect 364996 700806 365024 703520
rect 364984 700800 365036 700806
rect 364984 700742 365036 700748
rect 397472 700738 397500 703520
rect 397460 700732 397512 700738
rect 397460 700674 397512 700680
rect 413664 700670 413692 703520
rect 413652 700664 413704 700670
rect 413652 700606 413704 700612
rect 429856 700602 429884 703520
rect 429844 700596 429896 700602
rect 429844 700538 429896 700544
rect 462332 700534 462360 703520
rect 478524 702434 478552 703520
rect 477512 702406 478552 702434
rect 462320 700528 462372 700534
rect 462320 700470 462372 700476
rect 337658 376952 337714 376961
rect 337658 376887 337714 376896
rect 337672 376786 337700 376887
rect 337660 376780 337712 376786
rect 337660 376722 337712 376728
rect 337750 376000 337806 376009
rect 337750 375935 337806 375944
rect 337764 375426 337792 375935
rect 337752 375420 337804 375426
rect 337752 375362 337804 375368
rect 337474 373824 337530 373833
rect 337474 373759 337530 373768
rect 337488 372638 337516 373759
rect 337566 372872 337622 372881
rect 337566 372807 337622 372816
rect 337476 372632 337528 372638
rect 337476 372574 337528 372580
rect 337474 371104 337530 371113
rect 337474 371039 337530 371048
rect 337488 369986 337516 371039
rect 337476 369980 337528 369986
rect 337476 369922 337528 369928
rect 337474 368248 337530 368257
rect 337474 368183 337530 368192
rect 337488 367130 337516 368183
rect 337476 367124 337528 367130
rect 337476 367066 337528 367072
rect 337580 354674 337608 372807
rect 337750 370016 337806 370025
rect 337750 369951 337806 369960
rect 337764 369918 337792 369951
rect 337752 369912 337804 369918
rect 337752 369854 337804 369860
rect 337488 354646 337608 354674
rect 337382 348392 337438 348401
rect 337382 348327 337438 348336
rect 337396 338094 337424 348327
rect 337384 338088 337436 338094
rect 337384 338030 337436 338036
rect 299480 243772 299532 243778
rect 299480 243714 299532 243720
rect 294604 128308 294656 128314
rect 294604 128250 294656 128256
rect 291844 113076 291896 113082
rect 291844 113018 291896 113024
rect 337488 103494 337516 354646
rect 337750 350024 337806 350033
rect 337750 349959 337806 349968
rect 337764 349178 337792 349959
rect 337752 349172 337804 349178
rect 337752 349114 337804 349120
rect 337658 348120 337714 348129
rect 337658 348055 337714 348064
rect 337672 347818 337700 348055
rect 337660 347812 337712 347818
rect 337660 347754 337712 347760
rect 371238 338056 371294 338065
rect 371238 337991 371294 338000
rect 382370 338056 382426 338065
rect 382370 337991 382426 338000
rect 386418 338056 386474 338065
rect 386418 337991 386474 338000
rect 407118 338056 407174 338065
rect 407118 337991 407174 338000
rect 362958 337784 363014 337793
rect 362958 337719 363014 337728
rect 366362 337784 366418 337793
rect 366362 337719 366418 337728
rect 369858 337784 369914 337793
rect 369858 337719 369914 337728
rect 356058 337648 356114 337657
rect 356058 337583 356114 337592
rect 357438 337648 357494 337657
rect 357438 337583 357494 337592
rect 358818 337648 358874 337657
rect 358818 337583 358874 337592
rect 360198 337648 360254 337657
rect 360198 337583 360254 337592
rect 361578 337648 361634 337657
rect 361578 337583 361634 337592
rect 355324 337544 355376 337550
rect 355324 337486 355376 337492
rect 349804 337408 349856 337414
rect 349804 337350 349856 337356
rect 349816 245274 349844 337350
rect 352564 337340 352616 337346
rect 352564 337282 352616 337288
rect 351184 336796 351236 336802
rect 351184 336738 351236 336744
rect 349804 245268 349856 245274
rect 349804 245210 349856 245216
rect 341524 238808 341576 238814
rect 341524 238750 341576 238756
rect 341536 126954 341564 238750
rect 341524 126948 341576 126954
rect 341524 126890 341576 126896
rect 337476 103488 337528 103494
rect 337476 103430 337528 103436
rect 351196 67590 351224 336738
rect 351184 67584 351236 67590
rect 351184 67526 351236 67532
rect 352576 39234 352604 337282
rect 355336 243846 355364 337486
rect 355324 243840 355376 243846
rect 355324 243782 355376 243788
rect 356072 242350 356100 337583
rect 356060 242344 356112 242350
rect 356060 242286 356112 242292
rect 357452 238202 357480 337583
rect 357440 238196 357492 238202
rect 357440 238138 357492 238144
rect 358832 63510 358860 337583
rect 360212 78674 360240 337583
rect 361592 88330 361620 337583
rect 361580 88324 361632 88330
rect 361580 88266 361632 88272
rect 360200 78668 360252 78674
rect 360200 78610 360252 78616
rect 358820 63504 358872 63510
rect 358820 63446 358872 63452
rect 362972 52426 363000 337719
rect 363050 337648 363106 337657
rect 363050 337583 363106 337592
rect 365718 337648 365774 337657
rect 365718 337583 365774 337592
rect 363064 242282 363092 337583
rect 364984 337476 365036 337482
rect 364984 337418 365036 337424
rect 364522 336832 364578 336841
rect 364522 336767 364524 336776
rect 364576 336767 364578 336776
rect 364524 336738 364576 336744
rect 363052 242276 363104 242282
rect 363052 242218 363104 242224
rect 364996 238746 365024 337418
rect 365732 241126 365760 337583
rect 366376 242418 366404 337719
rect 369872 337686 369900 337719
rect 367744 337680 367796 337686
rect 367190 337648 367246 337657
rect 369860 337680 369912 337686
rect 367744 337622 367796 337628
rect 368478 337648 368534 337657
rect 367190 337583 367246 337592
rect 366364 242412 366416 242418
rect 366364 242354 366416 242360
rect 365720 241120 365772 241126
rect 365720 241062 365772 241068
rect 367204 241058 367232 337583
rect 367192 241052 367244 241058
rect 367192 240994 367244 241000
rect 364984 238740 365036 238746
rect 364984 238682 365036 238688
rect 367756 107642 367784 337622
rect 369860 337622 369912 337628
rect 369950 337648 370006 337657
rect 368478 337583 368534 337592
rect 369950 337583 370006 337592
rect 368492 240990 368520 337583
rect 369964 250714 369992 337583
rect 371252 337210 371280 337991
rect 375378 337920 375434 337929
rect 375378 337855 375434 337864
rect 379518 337920 379574 337929
rect 379518 337855 379520 337864
rect 372618 337784 372674 337793
rect 372618 337719 372674 337728
rect 371882 337648 371938 337657
rect 371882 337583 371938 337592
rect 371240 337204 371292 337210
rect 371240 337146 371292 337152
rect 371238 336832 371294 336841
rect 371238 336767 371294 336776
rect 371252 336122 371280 336767
rect 371240 336116 371292 336122
rect 371240 336058 371292 336064
rect 369952 250708 370004 250714
rect 369952 250650 370004 250656
rect 368480 240984 368532 240990
rect 368480 240926 368532 240932
rect 371896 143546 371924 337583
rect 372632 337550 372660 337719
rect 373998 337648 374054 337657
rect 373998 337583 374054 337592
rect 372620 337544 372672 337550
rect 372620 337486 372672 337492
rect 373264 336796 373316 336802
rect 373264 336738 373316 336744
rect 371884 143540 371936 143546
rect 371884 143482 371936 143488
rect 367744 107636 367796 107642
rect 367744 107578 367796 107584
rect 373276 93838 373304 336738
rect 374012 242486 374040 337583
rect 375392 337142 375420 337855
rect 379572 337855 379574 337864
rect 379520 337826 379572 337832
rect 378138 337784 378194 337793
rect 378138 337719 378194 337728
rect 380162 337784 380218 337793
rect 380162 337719 380218 337728
rect 375470 337648 375526 337657
rect 375470 337583 375526 337592
rect 376758 337648 376814 337657
rect 376758 337583 376814 337592
rect 375380 337136 375432 337142
rect 375380 337078 375432 337084
rect 375484 242554 375512 337583
rect 375472 242548 375524 242554
rect 375472 242490 375524 242496
rect 374000 242480 374052 242486
rect 374000 242422 374052 242428
rect 376772 242214 376800 337583
rect 376850 336832 376906 336841
rect 378152 336802 378180 337719
rect 379518 337104 379574 337113
rect 379440 337062 379518 337090
rect 379440 337006 379468 337062
rect 379518 337039 379574 337048
rect 379428 337000 379480 337006
rect 379428 336942 379480 336948
rect 379520 337000 379572 337006
rect 379520 336942 379572 336948
rect 376850 336767 376906 336776
rect 378140 336796 378192 336802
rect 376864 336598 376892 336767
rect 378140 336738 378192 336744
rect 376852 336592 376904 336598
rect 376852 336534 376904 336540
rect 379532 336462 379560 336942
rect 379520 336456 379572 336462
rect 379520 336398 379572 336404
rect 376760 242208 376812 242214
rect 376760 242150 376812 242156
rect 373264 93832 373316 93838
rect 373264 93774 373316 93780
rect 362960 52420 363012 52426
rect 362960 52362 363012 52368
rect 352564 39228 352616 39234
rect 352564 39170 352616 39176
rect 290464 38140 290516 38146
rect 290464 38082 290516 38088
rect 380176 38010 380204 337719
rect 380990 337648 381046 337657
rect 380990 337583 381046 337592
rect 381004 249082 381032 337583
rect 382278 337376 382334 337385
rect 382278 337311 382334 337320
rect 382292 337278 382320 337311
rect 382280 337272 382332 337278
rect 382280 337214 382332 337220
rect 381544 337136 381596 337142
rect 381544 337078 381596 337084
rect 380992 249076 381044 249082
rect 380992 249018 381044 249024
rect 381556 240922 381584 337078
rect 382384 336054 382412 337991
rect 384302 337648 384358 337657
rect 384302 337583 384358 337592
rect 382924 337204 382976 337210
rect 382924 337146 382976 337152
rect 382372 336048 382424 336054
rect 382372 335990 382424 335996
rect 382936 242690 382964 337146
rect 383750 336968 383806 336977
rect 383750 336903 383752 336912
rect 383804 336903 383806 336912
rect 383752 336874 383804 336880
rect 382924 242684 382976 242690
rect 382924 242626 382976 242632
rect 381544 240916 381596 240922
rect 381544 240858 381596 240864
rect 380164 38004 380216 38010
rect 380164 37946 380216 37952
rect 384316 37942 384344 337583
rect 385038 337512 385094 337521
rect 385038 337447 385094 337456
rect 385052 337414 385080 337447
rect 385040 337408 385092 337414
rect 385040 337350 385092 337356
rect 385684 337340 385736 337346
rect 385684 337282 385736 337288
rect 384948 336864 385000 336870
rect 384948 336806 385000 336812
rect 384960 336530 384988 336806
rect 384948 336524 385000 336530
rect 384948 336466 385000 336472
rect 385696 137970 385724 337282
rect 386432 337210 386460 337991
rect 394698 337920 394754 337929
rect 394698 337855 394754 337864
rect 397458 337920 397514 337929
rect 397458 337855 397514 337864
rect 394712 337822 394740 337855
rect 394700 337816 394752 337822
rect 389178 337784 389234 337793
rect 388444 337748 388496 337754
rect 389178 337719 389234 337728
rect 391938 337784 391994 337793
rect 394700 337758 394752 337764
rect 391938 337719 391940 337728
rect 388444 337690 388496 337696
rect 387064 337680 387116 337686
rect 387064 337622 387116 337628
rect 386510 337240 386566 337249
rect 386420 337204 386472 337210
rect 386510 337175 386566 337184
rect 386420 337146 386472 337152
rect 386524 337142 386552 337175
rect 386512 337136 386564 337142
rect 386512 337078 386564 337084
rect 387076 198694 387104 337622
rect 387798 337512 387854 337521
rect 387798 337447 387854 337456
rect 387812 337414 387840 337447
rect 387800 337408 387852 337414
rect 387800 337350 387852 337356
rect 387798 337104 387854 337113
rect 387798 337039 387854 337048
rect 387812 337006 387840 337039
rect 387800 337000 387852 337006
rect 387800 336942 387852 336948
rect 388456 208350 388484 337690
rect 389192 337686 389220 337719
rect 391992 337719 391994 337728
rect 391940 337690 391992 337696
rect 389180 337680 389232 337686
rect 389180 337622 389232 337628
rect 390558 337648 390614 337657
rect 390558 337583 390614 337592
rect 393410 337648 393466 337657
rect 393410 337583 393466 337592
rect 395342 337648 395398 337657
rect 395342 337583 395398 337592
rect 390572 337346 390600 337583
rect 390560 337340 390612 337346
rect 390560 337282 390612 337288
rect 392582 337104 392638 337113
rect 392582 337039 392638 337048
rect 390558 336832 390614 336841
rect 390558 336767 390614 336776
rect 391204 336796 391256 336802
rect 390572 336666 390600 336767
rect 391204 336738 391256 336744
rect 390560 336660 390612 336666
rect 390560 336602 390612 336608
rect 391216 242622 391244 336738
rect 391204 242616 391256 242622
rect 391204 242558 391256 242564
rect 388444 208344 388496 208350
rect 388444 208286 388496 208292
rect 387064 198688 387116 198694
rect 387064 198630 387116 198636
rect 385684 137964 385736 137970
rect 385684 137906 385736 137912
rect 392596 38486 392624 337039
rect 393318 336968 393374 336977
rect 393318 336903 393374 336912
rect 393332 336802 393360 336903
rect 393320 336796 393372 336802
rect 393320 336738 393372 336744
rect 393424 251870 393452 337583
rect 393412 251864 393464 251870
rect 393412 251806 393464 251812
rect 395356 38826 395384 337583
rect 397472 337482 397500 337855
rect 398102 337648 398158 337657
rect 398102 337583 398158 337592
rect 399574 337648 399630 337657
rect 399574 337583 399630 337592
rect 397460 337476 397512 337482
rect 397460 337418 397512 337424
rect 396078 336968 396134 336977
rect 396078 336903 396134 336912
rect 396092 336870 396120 336903
rect 396080 336864 396132 336870
rect 396080 336806 396132 336812
rect 397458 336832 397514 336841
rect 397458 336767 397514 336776
rect 397472 336258 397500 336767
rect 397460 336252 397512 336258
rect 397460 336194 397512 336200
rect 398116 242758 398144 337583
rect 399484 336864 399536 336870
rect 399484 336806 399536 336812
rect 398104 242752 398156 242758
rect 398104 242694 398156 242700
rect 399496 38962 399524 336806
rect 399588 269822 399616 337583
rect 405738 336968 405794 336977
rect 402244 336932 402296 336938
rect 407132 336938 407160 337991
rect 412638 337648 412694 337657
rect 412638 337583 412694 337592
rect 415398 337648 415454 337657
rect 415398 337583 415454 337592
rect 417422 337648 417478 337657
rect 417422 337583 417478 337592
rect 420918 337648 420974 337657
rect 420918 337583 420974 337592
rect 427818 337648 427874 337657
rect 427818 337583 427874 337592
rect 430578 337648 430634 337657
rect 430578 337583 430634 337592
rect 434718 337648 434774 337657
rect 434718 337583 434774 337592
rect 437478 337648 437534 337657
rect 437478 337583 437534 337592
rect 445758 337648 445814 337657
rect 445758 337583 445814 337592
rect 409878 337240 409934 337249
rect 409878 337175 409934 337184
rect 405738 336903 405794 336912
rect 407120 336932 407172 336938
rect 402244 336874 402296 336880
rect 399576 269816 399628 269822
rect 399576 269758 399628 269764
rect 399484 38956 399536 38962
rect 399484 38898 399536 38904
rect 402256 38894 402284 336874
rect 405752 336870 405780 336903
rect 407120 336874 407172 336880
rect 409144 336932 409196 336938
rect 409144 336874 409196 336880
rect 405740 336864 405792 336870
rect 403254 336832 403310 336841
rect 405740 336806 405792 336812
rect 406384 336864 406436 336870
rect 406384 336806 406436 336812
rect 403254 336767 403310 336776
rect 403268 336394 403296 336767
rect 403256 336388 403308 336394
rect 403256 336330 403308 336336
rect 406396 39098 406424 336806
rect 406384 39092 406436 39098
rect 406384 39034 406436 39040
rect 409156 39030 409184 336874
rect 409892 336326 409920 337175
rect 411904 337000 411956 337006
rect 411904 336942 411956 336948
rect 409880 336320 409932 336326
rect 409880 336262 409932 336268
rect 411916 39166 411944 336942
rect 412652 240854 412680 337583
rect 412640 240848 412692 240854
rect 412640 240790 412692 240796
rect 415412 185638 415440 337583
rect 417436 187678 417464 337583
rect 417424 187672 417476 187678
rect 417424 187614 417476 187620
rect 415400 185632 415452 185638
rect 415400 185574 415452 185580
rect 411904 39160 411956 39166
rect 411904 39102 411956 39108
rect 409144 39024 409196 39030
rect 409144 38966 409196 38972
rect 402244 38888 402296 38894
rect 402244 38830 402296 38836
rect 395344 38820 395396 38826
rect 395344 38762 395396 38768
rect 420932 38758 420960 337583
rect 422942 337376 422998 337385
rect 422942 337311 422998 337320
rect 422956 336870 422984 337311
rect 425058 336968 425114 336977
rect 425058 336903 425060 336912
rect 425112 336903 425114 336912
rect 425060 336874 425112 336880
rect 422944 336864 422996 336870
rect 422944 336806 422996 336812
rect 427832 204950 427860 337583
rect 430592 243710 430620 337583
rect 433338 337104 433394 337113
rect 433338 337039 433340 337048
rect 433392 337039 433394 337048
rect 433340 337010 433392 337016
rect 430580 243704 430632 243710
rect 430580 243646 430632 243652
rect 427820 204944 427872 204950
rect 427820 204886 427872 204892
rect 420920 38752 420972 38758
rect 420920 38694 420972 38700
rect 434732 38690 434760 337583
rect 437492 245138 437520 337583
rect 442998 337240 443054 337249
rect 442998 337175 443054 337184
rect 440238 337104 440294 337113
rect 440238 337039 440294 337048
rect 440252 337006 440280 337039
rect 440240 337000 440292 337006
rect 440240 336942 440292 336948
rect 443012 336190 443040 337175
rect 443000 336184 443052 336190
rect 443000 336126 443052 336132
rect 437480 245132 437532 245138
rect 437480 245074 437532 245080
rect 445772 243642 445800 337583
rect 477512 245070 477540 702406
rect 494808 700398 494836 703520
rect 527192 700466 527220 703520
rect 543476 702434 543504 703520
rect 542372 702406 543504 702434
rect 527180 700460 527232 700466
rect 527180 700402 527232 700408
rect 494796 700392 494848 700398
rect 494796 700334 494848 700340
rect 479524 456816 479576 456822
rect 479524 456758 479576 456764
rect 479536 247858 479564 456758
rect 486424 418192 486476 418198
rect 486424 418134 486476 418140
rect 482284 404388 482336 404394
rect 482284 404330 482336 404336
rect 480904 351960 480956 351966
rect 480904 351902 480956 351908
rect 479524 247852 479576 247858
rect 479524 247794 479576 247800
rect 480916 247722 480944 351902
rect 482296 247790 482324 404330
rect 483664 378208 483716 378214
rect 483664 378150 483716 378156
rect 483676 250578 483704 378150
rect 485044 364404 485096 364410
rect 485044 364346 485096 364352
rect 483664 250572 483716 250578
rect 483664 250514 483716 250520
rect 482284 247784 482336 247790
rect 482284 247726 482336 247732
rect 480904 247716 480956 247722
rect 480904 247658 480956 247664
rect 477500 245064 477552 245070
rect 477500 245006 477552 245012
rect 485056 245002 485084 364346
rect 486436 250646 486464 418134
rect 486424 250640 486476 250646
rect 486424 250582 486476 250588
rect 542372 250510 542400 702406
rect 559668 700330 559696 703520
rect 559656 700324 559708 700330
rect 559656 700266 559708 700272
rect 580170 697232 580226 697241
rect 580170 697167 580226 697176
rect 580184 696998 580212 697167
rect 580172 696992 580224 696998
rect 580172 696934 580224 696940
rect 580262 683904 580318 683913
rect 580262 683839 580318 683848
rect 580172 670744 580224 670750
rect 580170 670712 580172 670721
rect 580224 670712 580226 670721
rect 580170 670647 580226 670656
rect 580170 644056 580226 644065
rect 580170 643991 580226 644000
rect 580184 643142 580212 643991
rect 580172 643136 580224 643142
rect 580172 643078 580224 643084
rect 579986 630864 580042 630873
rect 579986 630799 580042 630808
rect 580000 630698 580028 630799
rect 579988 630692 580040 630698
rect 579988 630634 580040 630640
rect 580170 617536 580226 617545
rect 580170 617471 580226 617480
rect 580184 616894 580212 617471
rect 580172 616888 580224 616894
rect 580172 616830 580224 616836
rect 580170 591016 580226 591025
rect 580170 590951 580226 590960
rect 580184 590714 580212 590951
rect 580172 590708 580224 590714
rect 580172 590650 580224 590656
rect 579894 564360 579950 564369
rect 579894 564295 579950 564304
rect 579908 563106 579936 564295
rect 579896 563100 579948 563106
rect 579896 563042 579948 563048
rect 580170 537840 580226 537849
rect 580170 537775 580226 537784
rect 580184 536858 580212 537775
rect 580172 536852 580224 536858
rect 580172 536794 580224 536800
rect 580170 524512 580226 524521
rect 580170 524447 580172 524456
rect 580224 524447 580226 524456
rect 580172 524418 580224 524424
rect 580170 511320 580226 511329
rect 580170 511255 580226 511264
rect 580184 510678 580212 511255
rect 580172 510672 580224 510678
rect 580172 510614 580224 510620
rect 580170 484664 580226 484673
rect 580170 484599 580226 484608
rect 580184 484430 580212 484599
rect 580172 484424 580224 484430
rect 580172 484366 580224 484372
rect 579618 458144 579674 458153
rect 579618 458079 579674 458088
rect 579632 456822 579660 458079
rect 579620 456816 579672 456822
rect 579620 456758 579672 456764
rect 579710 418296 579766 418305
rect 579710 418231 579766 418240
rect 579724 418198 579752 418231
rect 579712 418192 579764 418198
rect 579712 418134 579764 418140
rect 580170 404968 580226 404977
rect 580170 404903 580226 404912
rect 580184 404394 580212 404903
rect 580172 404388 580224 404394
rect 580172 404330 580224 404336
rect 580170 378448 580226 378457
rect 580170 378383 580226 378392
rect 580184 378214 580212 378383
rect 580172 378208 580224 378214
rect 580172 378150 580224 378156
rect 580170 365120 580226 365129
rect 580170 365055 580226 365064
rect 580184 364410 580212 365055
rect 580172 364404 580224 364410
rect 580172 364346 580224 364352
rect 580172 351960 580224 351966
rect 580170 351928 580172 351937
rect 580224 351928 580226 351937
rect 580170 351863 580226 351872
rect 580276 338910 580304 683839
rect 580354 577688 580410 577697
rect 580354 577623 580410 577632
rect 580264 338904 580316 338910
rect 580264 338846 580316 338852
rect 580368 338842 580396 577623
rect 580538 471472 580594 471481
rect 580538 471407 580594 471416
rect 580446 431624 580502 431633
rect 580446 431559 580502 431568
rect 580356 338836 580408 338842
rect 580356 338778 580408 338784
rect 579986 325272 580042 325281
rect 579986 325207 580042 325216
rect 580000 324358 580028 325207
rect 579988 324352 580040 324358
rect 579988 324294 580040 324300
rect 580170 312080 580226 312089
rect 580170 312015 580226 312024
rect 580184 311914 580212 312015
rect 580172 311908 580224 311914
rect 580172 311850 580224 311856
rect 580170 298752 580226 298761
rect 580170 298687 580226 298696
rect 580184 298178 580212 298687
rect 580172 298172 580224 298178
rect 580172 298114 580224 298120
rect 580170 272232 580226 272241
rect 580170 272167 580226 272176
rect 580184 271930 580212 272167
rect 580172 271924 580224 271930
rect 580172 271866 580224 271872
rect 580170 258904 580226 258913
rect 580170 258839 580226 258848
rect 580184 258126 580212 258839
rect 580172 258120 580224 258126
rect 580172 258062 580224 258068
rect 542360 250504 542412 250510
rect 542360 250446 542412 250452
rect 579618 245576 579674 245585
rect 579618 245511 579674 245520
rect 485044 244996 485096 245002
rect 485044 244938 485096 244944
rect 445760 243636 445812 243642
rect 445760 243578 445812 243584
rect 579632 243574 579660 245511
rect 580460 244934 580488 431559
rect 580552 338774 580580 471407
rect 580540 338768 580592 338774
rect 580540 338710 580592 338716
rect 580448 244928 580500 244934
rect 580448 244870 580500 244876
rect 579620 243568 579672 243574
rect 579620 243510 579672 243516
rect 580172 240100 580224 240106
rect 580172 240042 580224 240048
rect 580184 229094 580212 240042
rect 580632 239760 580684 239766
rect 580632 239702 580684 239708
rect 580540 239692 580592 239698
rect 580540 239634 580592 239640
rect 580264 239556 580316 239562
rect 580264 239498 580316 239504
rect 580276 233866 580304 239498
rect 580448 239488 580500 239494
rect 580448 239430 580500 239436
rect 580356 239420 580408 239426
rect 580356 239362 580408 239368
rect 580368 235550 580396 239362
rect 580356 235544 580408 235550
rect 580356 235486 580408 235492
rect 580276 233838 580396 233866
rect 580184 229066 580304 229094
rect 579804 206984 579856 206990
rect 579804 206926 579856 206932
rect 579816 205737 579844 206926
rect 579802 205728 579858 205737
rect 579802 205663 579858 205672
rect 579620 193180 579672 193186
rect 579620 193122 579672 193128
rect 579632 192545 579660 193122
rect 579618 192536 579674 192545
rect 579618 192471 579674 192480
rect 580172 167000 580224 167006
rect 580172 166942 580224 166948
rect 580184 165889 580212 166942
rect 580170 165880 580226 165889
rect 580170 165815 580226 165824
rect 580172 139392 580224 139398
rect 580170 139360 580172 139369
rect 580224 139360 580226 139369
rect 580170 139295 580226 139304
rect 580172 126948 580224 126954
rect 580172 126890 580224 126896
rect 580184 126041 580212 126890
rect 580170 126032 580226 126041
rect 580170 125967 580226 125976
rect 579620 113144 579672 113150
rect 579620 113086 579672 113092
rect 579632 112849 579660 113086
rect 579618 112840 579674 112849
rect 579618 112775 579674 112784
rect 580172 100700 580224 100706
rect 580172 100642 580224 100648
rect 580184 99521 580212 100642
rect 580170 99512 580226 99521
rect 580170 99447 580226 99456
rect 579620 86964 579672 86970
rect 579620 86906 579672 86912
rect 579632 86193 579660 86906
rect 579618 86184 579674 86193
rect 579618 86119 579674 86128
rect 580172 73160 580224 73166
rect 580172 73102 580224 73108
rect 580184 73001 580212 73102
rect 580170 72992 580226 73001
rect 580170 72927 580226 72936
rect 580172 46912 580224 46918
rect 580172 46854 580224 46860
rect 580184 46345 580212 46854
rect 580170 46336 580226 46345
rect 580170 46271 580226 46280
rect 434720 38684 434772 38690
rect 434720 38626 434772 38632
rect 392584 38480 392636 38486
rect 392584 38422 392636 38428
rect 384304 37936 384356 37942
rect 384304 37878 384356 37884
rect 580170 33144 580226 33153
rect 273904 33108 273956 33114
rect 580170 33079 580172 33088
rect 273904 33050 273956 33056
rect 580224 33079 580226 33088
rect 580172 33050 580224 33056
rect 580276 19825 580304 229066
rect 580368 59673 580396 233838
rect 580460 152697 580488 239430
rect 580552 179217 580580 239634
rect 580644 219065 580672 239702
rect 580724 235544 580776 235550
rect 580724 235486 580776 235492
rect 580736 232393 580764 235486
rect 580722 232384 580778 232393
rect 580722 232319 580778 232328
rect 580630 219056 580686 219065
rect 580630 218991 580686 219000
rect 580538 179208 580594 179217
rect 580538 179143 580594 179152
rect 580446 152688 580502 152697
rect 580446 152623 580502 152632
rect 580354 59664 580410 59673
rect 580354 59599 580410 59608
rect 580262 19816 580318 19825
rect 580262 19751 580318 19760
rect 265624 6860 265676 6866
rect 265624 6802 265676 6808
rect 580172 6860 580224 6866
rect 580172 6802 580224 6808
rect 580184 6633 580212 6802
rect 580170 6624 580226 6633
rect 580170 6559 580226 6568
rect 582196 3596 582248 3602
rect 582196 3538 582248 3544
rect 183468 3528 183520 3534
rect 183468 3470 183520 3476
rect 173900 3460 173952 3466
rect 173900 3402 173952 3408
rect 180708 3460 180760 3466
rect 180708 3402 180760 3408
rect 581000 3460 581052 3466
rect 581000 3402 581052 3408
rect 124680 2848 124732 2854
rect 124680 2790 124732 2796
rect 128544 2848 128596 2854
rect 128544 2790 128596 2796
rect 124692 480 124720 2790
rect 581012 480 581040 3402
rect 582208 480 582236 3538
rect 583392 3528 583444 3534
rect 583392 3470 583444 3476
rect 583404 480 583432 3470
rect 542 -960 654 480
rect 1646 -960 1758 480
rect 2842 -960 2954 480
rect 4038 -960 4150 480
rect 5234 -960 5346 480
rect 6430 -960 6542 480
rect 7626 -960 7738 480
rect 8730 -960 8842 480
rect 9926 -960 10038 480
rect 11122 -960 11234 480
rect 12318 -960 12430 480
rect 13514 -960 13626 480
rect 14710 -960 14822 480
rect 15906 -960 16018 480
rect 17010 -960 17122 480
rect 18206 -960 18318 480
rect 19402 -960 19514 480
rect 20598 -960 20710 480
rect 21794 -960 21906 480
rect 22990 -960 23102 480
rect 24186 -960 24298 480
rect 25290 -960 25402 480
rect 26486 -960 26598 480
rect 27682 -960 27794 480
rect 28878 -960 28990 480
rect 30074 -960 30186 480
rect 31270 -960 31382 480
rect 32374 -960 32486 480
rect 33570 -960 33682 480
rect 34766 -960 34878 480
rect 35962 -960 36074 480
rect 37158 -960 37270 480
rect 38354 -960 38466 480
rect 39550 -960 39662 480
rect 40654 -960 40766 480
rect 41850 -960 41962 480
rect 43046 -960 43158 480
rect 44242 -960 44354 480
rect 45438 -960 45550 480
rect 46634 -960 46746 480
rect 47830 -960 47942 480
rect 48934 -960 49046 480
rect 50130 -960 50242 480
rect 51326 -960 51438 480
rect 52522 -960 52634 480
rect 53718 -960 53830 480
rect 54914 -960 55026 480
rect 56018 -960 56130 480
rect 57214 -960 57326 480
rect 58410 -960 58522 480
rect 59606 -960 59718 480
rect 60802 -960 60914 480
rect 61998 -960 62110 480
rect 63194 -960 63306 480
rect 64298 -960 64410 480
rect 65494 -960 65606 480
rect 66690 -960 66802 480
rect 67886 -960 67998 480
rect 69082 -960 69194 480
rect 70278 -960 70390 480
rect 71474 -960 71586 480
rect 72578 -960 72690 480
rect 73774 -960 73886 480
rect 74970 -960 75082 480
rect 76166 -960 76278 480
rect 77362 -960 77474 480
rect 78558 -960 78670 480
rect 79662 -960 79774 480
rect 80858 -960 80970 480
rect 82054 -960 82166 480
rect 83250 -960 83362 480
rect 84446 -960 84558 480
rect 85642 -960 85754 480
rect 86838 -960 86950 480
rect 87942 -960 88054 480
rect 89138 -960 89250 480
rect 90334 -960 90446 480
rect 91530 -960 91642 480
rect 92726 -960 92838 480
rect 93922 -960 94034 480
rect 95118 -960 95230 480
rect 96222 -960 96334 480
rect 97418 -960 97530 480
rect 98614 -960 98726 480
rect 99810 -960 99922 480
rect 101006 -960 101118 480
rect 102202 -960 102314 480
rect 103306 -960 103418 480
rect 104502 -960 104614 480
rect 105698 -960 105810 480
rect 106894 -960 107006 480
rect 108090 -960 108202 480
rect 109286 -960 109398 480
rect 110482 -960 110594 480
rect 111586 -960 111698 480
rect 112782 -960 112894 480
rect 113978 -960 114090 480
rect 115174 -960 115286 480
rect 116370 -960 116482 480
rect 117566 -960 117678 480
rect 118762 -960 118874 480
rect 119866 -960 119978 480
rect 121062 -960 121174 480
rect 122258 -960 122370 480
rect 123454 -960 123566 480
rect 124650 -960 124762 480
rect 125846 -960 125958 480
rect 126950 -960 127062 480
rect 128146 -960 128258 480
rect 129342 -960 129454 480
rect 130538 -960 130650 480
rect 131734 -960 131846 480
rect 132930 -960 133042 480
rect 134126 -960 134238 480
rect 135230 -960 135342 480
rect 136426 -960 136538 480
rect 137622 -960 137734 480
rect 138818 -960 138930 480
rect 140014 -960 140126 480
rect 141210 -960 141322 480
rect 142406 -960 142518 480
rect 143510 -960 143622 480
rect 144706 -960 144818 480
rect 145902 -960 146014 480
rect 147098 -960 147210 480
rect 148294 -960 148406 480
rect 149490 -960 149602 480
rect 150594 -960 150706 480
rect 151790 -960 151902 480
rect 152986 -960 153098 480
rect 154182 -960 154294 480
rect 155378 -960 155490 480
rect 156574 -960 156686 480
rect 157770 -960 157882 480
rect 158874 -960 158986 480
rect 160070 -960 160182 480
rect 161266 -960 161378 480
rect 162462 -960 162574 480
rect 163658 -960 163770 480
rect 164854 -960 164966 480
rect 166050 -960 166162 480
rect 167154 -960 167266 480
rect 168350 -960 168462 480
rect 169546 -960 169658 480
rect 170742 -960 170854 480
rect 171938 -960 172050 480
rect 173134 -960 173246 480
rect 174238 -960 174350 480
rect 175434 -960 175546 480
rect 176630 -960 176742 480
rect 177826 -960 177938 480
rect 179022 -960 179134 480
rect 180218 -960 180330 480
rect 181414 -960 181526 480
rect 182518 -960 182630 480
rect 183714 -960 183826 480
rect 184910 -960 185022 480
rect 186106 -960 186218 480
rect 187302 -960 187414 480
rect 188498 -960 188610 480
rect 189694 -960 189806 480
rect 190798 -960 190910 480
rect 191994 -960 192106 480
rect 193190 -960 193302 480
rect 194386 -960 194498 480
rect 195582 -960 195694 480
rect 196778 -960 196890 480
rect 197882 -960 197994 480
rect 199078 -960 199190 480
rect 200274 -960 200386 480
rect 201470 -960 201582 480
rect 202666 -960 202778 480
rect 203862 -960 203974 480
rect 205058 -960 205170 480
rect 206162 -960 206274 480
rect 207358 -960 207470 480
rect 208554 -960 208666 480
rect 209750 -960 209862 480
rect 210946 -960 211058 480
rect 212142 -960 212254 480
rect 213338 -960 213450 480
rect 214442 -960 214554 480
rect 215638 -960 215750 480
rect 216834 -960 216946 480
rect 218030 -960 218142 480
rect 219226 -960 219338 480
rect 220422 -960 220534 480
rect 221526 -960 221638 480
rect 222722 -960 222834 480
rect 223918 -960 224030 480
rect 225114 -960 225226 480
rect 226310 -960 226422 480
rect 227506 -960 227618 480
rect 228702 -960 228814 480
rect 229806 -960 229918 480
rect 231002 -960 231114 480
rect 232198 -960 232310 480
rect 233394 -960 233506 480
rect 234590 -960 234702 480
rect 235786 -960 235898 480
rect 236982 -960 237094 480
rect 238086 -960 238198 480
rect 239282 -960 239394 480
rect 240478 -960 240590 480
rect 241674 -960 241786 480
rect 242870 -960 242982 480
rect 244066 -960 244178 480
rect 245170 -960 245282 480
rect 246366 -960 246478 480
rect 247562 -960 247674 480
rect 248758 -960 248870 480
rect 249954 -960 250066 480
rect 251150 -960 251262 480
rect 252346 -960 252458 480
rect 253450 -960 253562 480
rect 254646 -960 254758 480
rect 255842 -960 255954 480
rect 257038 -960 257150 480
rect 258234 -960 258346 480
rect 259430 -960 259542 480
rect 260626 -960 260738 480
rect 261730 -960 261842 480
rect 262926 -960 263038 480
rect 264122 -960 264234 480
rect 265318 -960 265430 480
rect 266514 -960 266626 480
rect 267710 -960 267822 480
rect 268814 -960 268926 480
rect 270010 -960 270122 480
rect 271206 -960 271318 480
rect 272402 -960 272514 480
rect 273598 -960 273710 480
rect 274794 -960 274906 480
rect 275990 -960 276102 480
rect 277094 -960 277206 480
rect 278290 -960 278402 480
rect 279486 -960 279598 480
rect 280682 -960 280794 480
rect 281878 -960 281990 480
rect 283074 -960 283186 480
rect 284270 -960 284382 480
rect 285374 -960 285486 480
rect 286570 -960 286682 480
rect 287766 -960 287878 480
rect 288962 -960 289074 480
rect 290158 -960 290270 480
rect 291354 -960 291466 480
rect 292550 -960 292662 480
rect 293654 -960 293766 480
rect 294850 -960 294962 480
rect 296046 -960 296158 480
rect 297242 -960 297354 480
rect 298438 -960 298550 480
rect 299634 -960 299746 480
rect 300738 -960 300850 480
rect 301934 -960 302046 480
rect 303130 -960 303242 480
rect 304326 -960 304438 480
rect 305522 -960 305634 480
rect 306718 -960 306830 480
rect 307914 -960 308026 480
rect 309018 -960 309130 480
rect 310214 -960 310326 480
rect 311410 -960 311522 480
rect 312606 -960 312718 480
rect 313802 -960 313914 480
rect 314998 -960 315110 480
rect 316194 -960 316306 480
rect 317298 -960 317410 480
rect 318494 -960 318606 480
rect 319690 -960 319802 480
rect 320886 -960 320998 480
rect 322082 -960 322194 480
rect 323278 -960 323390 480
rect 324382 -960 324494 480
rect 325578 -960 325690 480
rect 326774 -960 326886 480
rect 327970 -960 328082 480
rect 329166 -960 329278 480
rect 330362 -960 330474 480
rect 331558 -960 331670 480
rect 332662 -960 332774 480
rect 333858 -960 333970 480
rect 335054 -960 335166 480
rect 336250 -960 336362 480
rect 337446 -960 337558 480
rect 338642 -960 338754 480
rect 339838 -960 339950 480
rect 340942 -960 341054 480
rect 342138 -960 342250 480
rect 343334 -960 343446 480
rect 344530 -960 344642 480
rect 345726 -960 345838 480
rect 346922 -960 347034 480
rect 348026 -960 348138 480
rect 349222 -960 349334 480
rect 350418 -960 350530 480
rect 351614 -960 351726 480
rect 352810 -960 352922 480
rect 354006 -960 354118 480
rect 355202 -960 355314 480
rect 356306 -960 356418 480
rect 357502 -960 357614 480
rect 358698 -960 358810 480
rect 359894 -960 360006 480
rect 361090 -960 361202 480
rect 362286 -960 362398 480
rect 363482 -960 363594 480
rect 364586 -960 364698 480
rect 365782 -960 365894 480
rect 366978 -960 367090 480
rect 368174 -960 368286 480
rect 369370 -960 369482 480
rect 370566 -960 370678 480
rect 371670 -960 371782 480
rect 372866 -960 372978 480
rect 374062 -960 374174 480
rect 375258 -960 375370 480
rect 376454 -960 376566 480
rect 377650 -960 377762 480
rect 378846 -960 378958 480
rect 379950 -960 380062 480
rect 381146 -960 381258 480
rect 382342 -960 382454 480
rect 383538 -960 383650 480
rect 384734 -960 384846 480
rect 385930 -960 386042 480
rect 387126 -960 387238 480
rect 388230 -960 388342 480
rect 389426 -960 389538 480
rect 390622 -960 390734 480
rect 391818 -960 391930 480
rect 393014 -960 393126 480
rect 394210 -960 394322 480
rect 395314 -960 395426 480
rect 396510 -960 396622 480
rect 397706 -960 397818 480
rect 398902 -960 399014 480
rect 400098 -960 400210 480
rect 401294 -960 401406 480
rect 402490 -960 402602 480
rect 403594 -960 403706 480
rect 404790 -960 404902 480
rect 405986 -960 406098 480
rect 407182 -960 407294 480
rect 408378 -960 408490 480
rect 409574 -960 409686 480
rect 410770 -960 410882 480
rect 411874 -960 411986 480
rect 413070 -960 413182 480
rect 414266 -960 414378 480
rect 415462 -960 415574 480
rect 416658 -960 416770 480
rect 417854 -960 417966 480
rect 418958 -960 419070 480
rect 420154 -960 420266 480
rect 421350 -960 421462 480
rect 422546 -960 422658 480
rect 423742 -960 423854 480
rect 424938 -960 425050 480
rect 426134 -960 426246 480
rect 427238 -960 427350 480
rect 428434 -960 428546 480
rect 429630 -960 429742 480
rect 430826 -960 430938 480
rect 432022 -960 432134 480
rect 433218 -960 433330 480
rect 434414 -960 434526 480
rect 435518 -960 435630 480
rect 436714 -960 436826 480
rect 437910 -960 438022 480
rect 439106 -960 439218 480
rect 440302 -960 440414 480
rect 441498 -960 441610 480
rect 442602 -960 442714 480
rect 443798 -960 443910 480
rect 444994 -960 445106 480
rect 446190 -960 446302 480
rect 447386 -960 447498 480
rect 448582 -960 448694 480
rect 449778 -960 449890 480
rect 450882 -960 450994 480
rect 452078 -960 452190 480
rect 453274 -960 453386 480
rect 454470 -960 454582 480
rect 455666 -960 455778 480
rect 456862 -960 456974 480
rect 458058 -960 458170 480
rect 459162 -960 459274 480
rect 460358 -960 460470 480
rect 461554 -960 461666 480
rect 462750 -960 462862 480
rect 463946 -960 464058 480
rect 465142 -960 465254 480
rect 466246 -960 466358 480
rect 467442 -960 467554 480
rect 468638 -960 468750 480
rect 469834 -960 469946 480
rect 471030 -960 471142 480
rect 472226 -960 472338 480
rect 473422 -960 473534 480
rect 474526 -960 474638 480
rect 475722 -960 475834 480
rect 476918 -960 477030 480
rect 478114 -960 478226 480
rect 479310 -960 479422 480
rect 480506 -960 480618 480
rect 481702 -960 481814 480
rect 482806 -960 482918 480
rect 484002 -960 484114 480
rect 485198 -960 485310 480
rect 486394 -960 486506 480
rect 487590 -960 487702 480
rect 488786 -960 488898 480
rect 489890 -960 490002 480
rect 491086 -960 491198 480
rect 492282 -960 492394 480
rect 493478 -960 493590 480
rect 494674 -960 494786 480
rect 495870 -960 495982 480
rect 497066 -960 497178 480
rect 498170 -960 498282 480
rect 499366 -960 499478 480
rect 500562 -960 500674 480
rect 501758 -960 501870 480
rect 502954 -960 503066 480
rect 504150 -960 504262 480
rect 505346 -960 505458 480
rect 506450 -960 506562 480
rect 507646 -960 507758 480
rect 508842 -960 508954 480
rect 510038 -960 510150 480
rect 511234 -960 511346 480
rect 512430 -960 512542 480
rect 513534 -960 513646 480
rect 514730 -960 514842 480
rect 515926 -960 516038 480
rect 517122 -960 517234 480
rect 518318 -960 518430 480
rect 519514 -960 519626 480
rect 520710 -960 520822 480
rect 521814 -960 521926 480
rect 523010 -960 523122 480
rect 524206 -960 524318 480
rect 525402 -960 525514 480
rect 526598 -960 526710 480
rect 527794 -960 527906 480
rect 528990 -960 529102 480
rect 530094 -960 530206 480
rect 531290 -960 531402 480
rect 532486 -960 532598 480
rect 533682 -960 533794 480
rect 534878 -960 534990 480
rect 536074 -960 536186 480
rect 537178 -960 537290 480
rect 538374 -960 538486 480
rect 539570 -960 539682 480
rect 540766 -960 540878 480
rect 541962 -960 542074 480
rect 543158 -960 543270 480
rect 544354 -960 544466 480
rect 545458 -960 545570 480
rect 546654 -960 546766 480
rect 547850 -960 547962 480
rect 549046 -960 549158 480
rect 550242 -960 550354 480
rect 551438 -960 551550 480
rect 552634 -960 552746 480
rect 553738 -960 553850 480
rect 554934 -960 555046 480
rect 556130 -960 556242 480
rect 557326 -960 557438 480
rect 558522 -960 558634 480
rect 559718 -960 559830 480
rect 560822 -960 560934 480
rect 562018 -960 562130 480
rect 563214 -960 563326 480
rect 564410 -960 564522 480
rect 565606 -960 565718 480
rect 566802 -960 566914 480
rect 567998 -960 568110 480
rect 569102 -960 569214 480
rect 570298 -960 570410 480
rect 571494 -960 571606 480
rect 572690 -960 572802 480
rect 573886 -960 573998 480
rect 575082 -960 575194 480
rect 576278 -960 576390 480
rect 577382 -960 577494 480
rect 578578 -960 578690 480
rect 579774 -960 579886 480
rect 580970 -960 581082 480
rect 582166 -960 582278 480
rect 583362 -960 583474 480
<< via2 >>
rect 2778 684256 2834 684312
rect 3422 671200 3478 671256
rect 3330 606056 3386 606112
rect 3330 579944 3386 580000
rect 3330 553832 3386 553888
rect 3330 527856 3386 527912
rect 3330 514820 3386 514856
rect 3330 514800 3332 514820
rect 3332 514800 3384 514820
rect 3384 514800 3386 514820
rect 2870 501744 2926 501800
rect 3330 475632 3386 475688
rect 3330 462576 3386 462632
rect 3330 449520 3386 449576
rect 3146 423544 3202 423600
rect 3330 397468 3332 397488
rect 3332 397468 3384 397488
rect 3384 397468 3386 397488
rect 3330 397432 3386 397468
rect 3330 371320 3386 371376
rect 3054 345344 3110 345400
rect 3514 658144 3570 658200
rect 3514 632068 3516 632088
rect 3516 632068 3568 632088
rect 3568 632068 3570 632088
rect 3514 632032 3570 632068
rect 3514 619112 3570 619168
rect 3606 566888 3662 566944
rect 3698 410488 3754 410544
rect 3422 319232 3478 319288
rect 3422 306176 3478 306232
rect 3422 293120 3478 293176
rect 3054 267144 3110 267200
rect 3422 254088 3478 254144
rect 3790 358400 3846 358456
rect 38382 376896 38438 376952
rect 37554 375944 37610 376000
rect 3422 241032 3478 241088
rect 3330 214920 3386 214976
rect 3054 201864 3110 201920
rect 3238 162832 3294 162888
rect 3146 110608 3202 110664
rect 3514 188844 3516 188864
rect 3516 188844 3568 188864
rect 3568 188844 3570 188864
rect 3514 188808 3570 188844
rect 3514 149776 3570 149832
rect 3514 136720 3570 136776
rect 3422 97552 3478 97608
rect 3146 84632 3202 84688
rect 3146 71612 3148 71632
rect 3148 71612 3200 71632
rect 3200 71612 3202 71632
rect 3146 71576 3202 71612
rect 3054 58520 3110 58576
rect 3422 45500 3424 45520
rect 3424 45500 3476 45520
rect 3476 45500 3478 45520
rect 3422 45464 3478 45500
rect 2870 32408 2926 32464
rect 3422 19352 3478 19408
rect 3422 6432 3478 6488
rect 36542 215736 36598 215792
rect 36634 210432 36690 210488
rect 36818 183368 36874 183424
rect 36726 177928 36782 177984
rect 36910 161608 36966 161664
rect 37094 145424 37150 145480
rect 37922 371048 37978 371104
rect 38198 349968 38254 350024
rect 37646 348064 37702 348120
rect 38750 373768 38806 373824
rect 38474 372816 38530 372872
rect 37738 199552 37794 199608
rect 37830 188672 37886 188728
rect 37738 150864 37794 150920
rect 37554 129104 37610 129160
rect 37922 167048 37978 167104
rect 38014 156304 38070 156360
rect 38014 134544 38070 134600
rect 38014 123800 38070 123856
rect 38106 112920 38162 112976
rect 38014 107480 38070 107536
rect 37830 102040 37886 102096
rect 37186 85856 37242 85912
rect 38014 74976 38070 75032
rect 38290 96736 38346 96792
rect 38382 80416 38438 80472
rect 38198 64232 38254 64288
rect 37002 53352 37058 53408
rect 38014 42608 38070 42664
rect 38658 369960 38714 370016
rect 38566 348336 38622 348392
rect 38842 368192 38898 368248
rect 38566 232056 38622 232112
rect 38566 69672 38622 69728
rect 38750 172488 38806 172544
rect 39210 204992 39266 205048
rect 39118 194112 39174 194168
rect 39026 139984 39082 140040
rect 38934 118360 38990 118416
rect 38842 91296 38898 91352
rect 38658 58792 38714 58848
rect 38566 45464 38622 45520
rect 77206 338000 77262 338056
rect 81254 338000 81310 338056
rect 59358 337864 59414 337920
rect 40406 337320 40462 337376
rect 40130 238040 40186 238096
rect 39486 226616 39542 226672
rect 39394 221176 39450 221232
rect 40590 242936 40646 242992
rect 43074 241576 43130 241632
rect 56506 337728 56562 337784
rect 57886 337728 57942 337784
rect 57978 337456 58034 337512
rect 60646 337728 60702 337784
rect 62118 337728 62174 337784
rect 64786 337728 64842 337784
rect 68834 337728 68890 337784
rect 69662 337728 69718 337784
rect 60002 337456 60058 337512
rect 60002 337184 60058 337240
rect 60738 337184 60794 337240
rect 45926 239808 45982 239864
rect 66166 337184 66222 337240
rect 67546 337184 67602 337240
rect 68926 337592 68982 337648
rect 78586 337864 78642 337920
rect 71318 337592 71374 337648
rect 74630 337592 74686 337648
rect 69662 336912 69718 336968
rect 70306 336796 70362 336832
rect 70306 336776 70308 336796
rect 70308 336776 70360 336796
rect 70360 336776 70362 336796
rect 75918 336776 75974 336832
rect 79966 337592 80022 337648
rect 82174 337592 82230 337648
rect 81346 337456 81402 337512
rect 84014 338000 84070 338056
rect 82910 337592 82966 337648
rect 73434 239808 73490 239864
rect 86866 337728 86922 337784
rect 87142 337728 87198 337784
rect 85486 337592 85542 337648
rect 85670 337592 85726 337648
rect 87050 337592 87106 337648
rect 50986 239672 51042 239728
rect 57702 239708 57704 239728
rect 57704 239708 57756 239728
rect 57756 239708 57758 239728
rect 57702 239672 57758 239708
rect 59174 239708 59176 239728
rect 59176 239708 59228 239728
rect 59228 239708 59230 239728
rect 59174 239672 59230 239708
rect 75826 239708 75828 239728
rect 75828 239708 75880 239728
rect 75880 239708 75882 239728
rect 75826 239672 75882 239708
rect 91006 338000 91062 338056
rect 89626 337728 89682 337784
rect 89718 337592 89774 337648
rect 93582 337864 93638 337920
rect 92386 337728 92442 337784
rect 91190 337592 91246 337648
rect 96618 337728 96674 337784
rect 93674 337592 93730 337648
rect 96342 337592 96398 337648
rect 95146 336796 95202 336832
rect 95146 336776 95148 336796
rect 95148 336776 95200 336796
rect 95200 336776 95202 336796
rect 96526 336776 96582 336832
rect 97998 338000 98054 338056
rect 99102 337592 99158 337648
rect 99286 337592 99342 337648
rect 104806 337728 104862 337784
rect 113178 337728 113234 337784
rect 117226 337728 117282 337784
rect 118606 337728 118662 337784
rect 102046 337592 102102 337648
rect 104898 337592 104954 337648
rect 108946 337592 109002 337648
rect 121274 336776 121330 336832
rect 122838 337728 122894 337784
rect 125598 337728 125654 337784
rect 131026 338000 131082 338056
rect 129646 336776 129702 336832
rect 133786 337728 133842 337784
rect 136546 337728 136602 337784
rect 139306 337728 139362 337784
rect 142066 337048 142122 337104
rect 143446 337728 143502 337784
rect 146206 337728 146262 337784
rect 168470 241576 168526 241632
rect 87142 239672 87198 239728
rect 237562 41112 237618 41168
rect 237746 40976 237802 41032
rect 237654 40840 237710 40896
rect 237930 57840 237986 57896
rect 237930 40840 237986 40896
rect 58254 39908 58310 39944
rect 58254 39888 58256 39908
rect 58256 39888 58308 39908
rect 58308 39888 58310 39908
rect 203338 38528 203394 38584
rect 207294 38392 207350 38448
rect 204718 38256 204774 38312
rect 200762 38120 200818 38176
rect 192850 37984 192906 38040
rect 188894 37848 188950 37904
rect 187606 37712 187662 37768
rect 215206 38528 215262 38584
rect 216494 38392 216550 38448
rect 238114 162288 238170 162344
rect 238758 122576 238814 122632
rect 238206 41112 238262 41168
rect 238114 40976 238170 41032
rect 238942 42472 238998 42528
rect 240138 227704 240194 227760
rect 239494 217640 239550 217696
rect 240138 177656 240194 177712
rect 239310 167592 239366 167648
rect 239218 147600 239274 147656
rect 239126 97552 239182 97608
rect 240322 82456 240378 82512
rect 240598 232736 240654 232792
rect 240598 192616 240654 192672
rect 240506 152632 240562 152688
rect 241150 237768 241206 237824
rect 240874 222672 240930 222728
rect 241242 212744 241298 212800
rect 241426 207712 241482 207768
rect 241426 202680 241482 202736
rect 241426 197648 241482 197704
rect 241426 187620 241428 187640
rect 241428 187620 241480 187640
rect 241480 187620 241482 187640
rect 241426 187584 241482 187620
rect 241426 182688 241482 182744
rect 241242 172624 241298 172680
rect 241058 157528 241114 157584
rect 241150 142568 241206 142624
rect 241426 137536 241482 137592
rect 240690 132504 240746 132560
rect 241426 127608 241482 127664
rect 240874 112512 240930 112568
rect 241426 107480 241482 107536
rect 241242 102448 241298 102504
rect 241426 92520 241482 92576
rect 241426 87488 241482 87544
rect 241242 77424 241298 77480
rect 240414 72392 240470 72448
rect 241426 67532 241428 67552
rect 241428 67532 241480 67552
rect 241480 67532 241482 67552
rect 241426 67496 241482 67532
rect 241242 62464 241298 62520
rect 241426 52420 241482 52456
rect 241426 52400 241428 52420
rect 241428 52400 241480 52420
rect 241480 52400 241482 52420
rect 240230 47368 240286 47424
rect 241702 117544 241758 117600
rect 265622 242936 265678 242992
rect 276662 238856 276718 238912
rect 283562 238720 283618 238776
rect 337658 376896 337714 376952
rect 337750 375944 337806 376000
rect 337474 373768 337530 373824
rect 337566 372816 337622 372872
rect 337474 371048 337530 371104
rect 337474 368192 337530 368248
rect 337750 369960 337806 370016
rect 337382 348336 337438 348392
rect 337750 349968 337806 350024
rect 337658 348064 337714 348120
rect 371238 338000 371294 338056
rect 382370 338000 382426 338056
rect 386418 338000 386474 338056
rect 407118 338000 407174 338056
rect 362958 337728 363014 337784
rect 366362 337728 366418 337784
rect 369858 337728 369914 337784
rect 356058 337592 356114 337648
rect 357438 337592 357494 337648
rect 358818 337592 358874 337648
rect 360198 337592 360254 337648
rect 361578 337592 361634 337648
rect 363050 337592 363106 337648
rect 365718 337592 365774 337648
rect 364522 336796 364578 336832
rect 364522 336776 364524 336796
rect 364524 336776 364576 336796
rect 364576 336776 364578 336796
rect 367190 337592 367246 337648
rect 368478 337592 368534 337648
rect 369950 337592 370006 337648
rect 375378 337864 375434 337920
rect 379518 337884 379574 337920
rect 379518 337864 379520 337884
rect 379520 337864 379572 337884
rect 379572 337864 379574 337884
rect 372618 337728 372674 337784
rect 371882 337592 371938 337648
rect 371238 336776 371294 336832
rect 373998 337592 374054 337648
rect 378138 337728 378194 337784
rect 380162 337728 380218 337784
rect 375470 337592 375526 337648
rect 376758 337592 376814 337648
rect 376850 336776 376906 336832
rect 379518 337048 379574 337104
rect 380990 337592 381046 337648
rect 382278 337320 382334 337376
rect 384302 337592 384358 337648
rect 383750 336932 383806 336968
rect 383750 336912 383752 336932
rect 383752 336912 383804 336932
rect 383804 336912 383806 336932
rect 385038 337456 385094 337512
rect 394698 337864 394754 337920
rect 397458 337864 397514 337920
rect 389178 337728 389234 337784
rect 391938 337748 391994 337784
rect 391938 337728 391940 337748
rect 391940 337728 391992 337748
rect 391992 337728 391994 337748
rect 386510 337184 386566 337240
rect 387798 337456 387854 337512
rect 387798 337048 387854 337104
rect 390558 337592 390614 337648
rect 393410 337592 393466 337648
rect 395342 337592 395398 337648
rect 392582 337048 392638 337104
rect 390558 336776 390614 336832
rect 393318 336912 393374 336968
rect 398102 337592 398158 337648
rect 399574 337592 399630 337648
rect 396078 336912 396134 336968
rect 397458 336776 397514 336832
rect 405738 336912 405794 336968
rect 412638 337592 412694 337648
rect 415398 337592 415454 337648
rect 417422 337592 417478 337648
rect 420918 337592 420974 337648
rect 427818 337592 427874 337648
rect 430578 337592 430634 337648
rect 434718 337592 434774 337648
rect 437478 337592 437534 337648
rect 445758 337592 445814 337648
rect 409878 337184 409934 337240
rect 403254 336776 403310 336832
rect 422942 337320 422998 337376
rect 425058 336932 425114 336968
rect 425058 336912 425060 336932
rect 425060 336912 425112 336932
rect 425112 336912 425114 336932
rect 433338 337068 433394 337104
rect 433338 337048 433340 337068
rect 433340 337048 433392 337068
rect 433392 337048 433394 337068
rect 442998 337184 443054 337240
rect 440238 337048 440294 337104
rect 580170 697176 580226 697232
rect 580262 683848 580318 683904
rect 580170 670692 580172 670712
rect 580172 670692 580224 670712
rect 580224 670692 580226 670712
rect 580170 670656 580226 670692
rect 580170 644000 580226 644056
rect 579986 630808 580042 630864
rect 580170 617480 580226 617536
rect 580170 590960 580226 591016
rect 579894 564304 579950 564360
rect 580170 537784 580226 537840
rect 580170 524476 580226 524512
rect 580170 524456 580172 524476
rect 580172 524456 580224 524476
rect 580224 524456 580226 524476
rect 580170 511264 580226 511320
rect 580170 484608 580226 484664
rect 579618 458088 579674 458144
rect 579710 418240 579766 418296
rect 580170 404912 580226 404968
rect 580170 378392 580226 378448
rect 580170 365064 580226 365120
rect 580170 351908 580172 351928
rect 580172 351908 580224 351928
rect 580224 351908 580226 351928
rect 580170 351872 580226 351908
rect 580354 577632 580410 577688
rect 580538 471416 580594 471472
rect 580446 431568 580502 431624
rect 579986 325216 580042 325272
rect 580170 312024 580226 312080
rect 580170 298696 580226 298752
rect 580170 272176 580226 272232
rect 580170 258848 580226 258904
rect 579618 245520 579674 245576
rect 579802 205672 579858 205728
rect 579618 192480 579674 192536
rect 580170 165824 580226 165880
rect 580170 139340 580172 139360
rect 580172 139340 580224 139360
rect 580224 139340 580226 139360
rect 580170 139304 580226 139340
rect 580170 125976 580226 126032
rect 579618 112784 579674 112840
rect 580170 99456 580226 99512
rect 579618 86128 579674 86184
rect 580170 72936 580226 72992
rect 580170 46280 580226 46336
rect 580170 33108 580226 33144
rect 580170 33088 580172 33108
rect 580172 33088 580224 33108
rect 580224 33088 580226 33108
rect 580722 232328 580778 232384
rect 580630 219000 580686 219056
rect 580538 179152 580594 179208
rect 580446 152632 580502 152688
rect 580354 59608 580410 59664
rect 580262 19760 580318 19816
rect 580170 6568 580226 6624
<< metal3 >>
rect -960 697220 480 697460
rect 580165 697234 580231 697237
rect 583520 697234 584960 697324
rect 580165 697232 584960 697234
rect 580165 697176 580170 697232
rect 580226 697176 584960 697232
rect 580165 697174 584960 697176
rect 580165 697171 580231 697174
rect 583520 697084 584960 697174
rect -960 684314 480 684404
rect 2773 684314 2839 684317
rect -960 684312 2839 684314
rect -960 684256 2778 684312
rect 2834 684256 2839 684312
rect -960 684254 2839 684256
rect -960 684164 480 684254
rect 2773 684251 2839 684254
rect 580257 683906 580323 683909
rect 583520 683906 584960 683996
rect 580257 683904 584960 683906
rect 580257 683848 580262 683904
rect 580318 683848 584960 683904
rect 580257 683846 584960 683848
rect 580257 683843 580323 683846
rect 583520 683756 584960 683846
rect -960 671258 480 671348
rect 3417 671258 3483 671261
rect -960 671256 3483 671258
rect -960 671200 3422 671256
rect 3478 671200 3483 671256
rect -960 671198 3483 671200
rect -960 671108 480 671198
rect 3417 671195 3483 671198
rect 580165 670714 580231 670717
rect 583520 670714 584960 670804
rect 580165 670712 584960 670714
rect 580165 670656 580170 670712
rect 580226 670656 584960 670712
rect 580165 670654 584960 670656
rect 580165 670651 580231 670654
rect 583520 670564 584960 670654
rect -960 658202 480 658292
rect 3509 658202 3575 658205
rect -960 658200 3575 658202
rect -960 658144 3514 658200
rect 3570 658144 3575 658200
rect -960 658142 3575 658144
rect -960 658052 480 658142
rect 3509 658139 3575 658142
rect 583520 657236 584960 657476
rect -960 644996 480 645236
rect 580165 644058 580231 644061
rect 583520 644058 584960 644148
rect 580165 644056 584960 644058
rect 580165 644000 580170 644056
rect 580226 644000 584960 644056
rect 580165 643998 584960 644000
rect 580165 643995 580231 643998
rect 583520 643908 584960 643998
rect -960 632090 480 632180
rect 3509 632090 3575 632093
rect -960 632088 3575 632090
rect -960 632032 3514 632088
rect 3570 632032 3575 632088
rect -960 632030 3575 632032
rect -960 631940 480 632030
rect 3509 632027 3575 632030
rect 579981 630866 580047 630869
rect 583520 630866 584960 630956
rect 579981 630864 584960 630866
rect 579981 630808 579986 630864
rect 580042 630808 584960 630864
rect 579981 630806 584960 630808
rect 579981 630803 580047 630806
rect 583520 630716 584960 630806
rect -960 619170 480 619260
rect 3509 619170 3575 619173
rect -960 619168 3575 619170
rect -960 619112 3514 619168
rect 3570 619112 3575 619168
rect -960 619110 3575 619112
rect -960 619020 480 619110
rect 3509 619107 3575 619110
rect 580165 617538 580231 617541
rect 583520 617538 584960 617628
rect 580165 617536 584960 617538
rect 580165 617480 580170 617536
rect 580226 617480 584960 617536
rect 580165 617478 584960 617480
rect 580165 617475 580231 617478
rect 583520 617388 584960 617478
rect -960 606114 480 606204
rect 3325 606114 3391 606117
rect -960 606112 3391 606114
rect -960 606056 3330 606112
rect 3386 606056 3391 606112
rect -960 606054 3391 606056
rect -960 605964 480 606054
rect 3325 606051 3391 606054
rect 583520 604060 584960 604300
rect -960 592908 480 593148
rect 580165 591018 580231 591021
rect 583520 591018 584960 591108
rect 580165 591016 584960 591018
rect 580165 590960 580170 591016
rect 580226 590960 584960 591016
rect 580165 590958 584960 590960
rect 580165 590955 580231 590958
rect 583520 590868 584960 590958
rect -960 580002 480 580092
rect 3325 580002 3391 580005
rect -960 580000 3391 580002
rect -960 579944 3330 580000
rect 3386 579944 3391 580000
rect -960 579942 3391 579944
rect -960 579852 480 579942
rect 3325 579939 3391 579942
rect 580349 577690 580415 577693
rect 583520 577690 584960 577780
rect 580349 577688 584960 577690
rect 580349 577632 580354 577688
rect 580410 577632 584960 577688
rect 580349 577630 584960 577632
rect 580349 577627 580415 577630
rect 583520 577540 584960 577630
rect -960 566946 480 567036
rect 3601 566946 3667 566949
rect -960 566944 3667 566946
rect -960 566888 3606 566944
rect 3662 566888 3667 566944
rect -960 566886 3667 566888
rect -960 566796 480 566886
rect 3601 566883 3667 566886
rect 579889 564362 579955 564365
rect 583520 564362 584960 564452
rect 579889 564360 584960 564362
rect 579889 564304 579894 564360
rect 579950 564304 584960 564360
rect 579889 564302 584960 564304
rect 579889 564299 579955 564302
rect 583520 564212 584960 564302
rect -960 553890 480 553980
rect 3325 553890 3391 553893
rect -960 553888 3391 553890
rect -960 553832 3330 553888
rect 3386 553832 3391 553888
rect -960 553830 3391 553832
rect -960 553740 480 553830
rect 3325 553827 3391 553830
rect 583520 551020 584960 551260
rect -960 540684 480 540924
rect 580165 537842 580231 537845
rect 583520 537842 584960 537932
rect 580165 537840 584960 537842
rect 580165 537784 580170 537840
rect 580226 537784 584960 537840
rect 580165 537782 584960 537784
rect 580165 537779 580231 537782
rect 583520 537692 584960 537782
rect -960 527914 480 528004
rect 3325 527914 3391 527917
rect -960 527912 3391 527914
rect -960 527856 3330 527912
rect 3386 527856 3391 527912
rect -960 527854 3391 527856
rect -960 527764 480 527854
rect 3325 527851 3391 527854
rect 580165 524514 580231 524517
rect 583520 524514 584960 524604
rect 580165 524512 584960 524514
rect 580165 524456 580170 524512
rect 580226 524456 584960 524512
rect 580165 524454 584960 524456
rect 580165 524451 580231 524454
rect 583520 524364 584960 524454
rect -960 514858 480 514948
rect 3325 514858 3391 514861
rect -960 514856 3391 514858
rect -960 514800 3330 514856
rect 3386 514800 3391 514856
rect -960 514798 3391 514800
rect -960 514708 480 514798
rect 3325 514795 3391 514798
rect 580165 511322 580231 511325
rect 583520 511322 584960 511412
rect 580165 511320 584960 511322
rect 580165 511264 580170 511320
rect 580226 511264 584960 511320
rect 580165 511262 584960 511264
rect 580165 511259 580231 511262
rect 583520 511172 584960 511262
rect -960 501802 480 501892
rect 2865 501802 2931 501805
rect -960 501800 2931 501802
rect -960 501744 2870 501800
rect 2926 501744 2931 501800
rect -960 501742 2931 501744
rect -960 501652 480 501742
rect 2865 501739 2931 501742
rect 583520 497844 584960 498084
rect -960 488596 480 488836
rect 580165 484666 580231 484669
rect 583520 484666 584960 484756
rect 580165 484664 584960 484666
rect 580165 484608 580170 484664
rect 580226 484608 584960 484664
rect 580165 484606 584960 484608
rect 580165 484603 580231 484606
rect 583520 484516 584960 484606
rect -960 475690 480 475780
rect 3325 475690 3391 475693
rect -960 475688 3391 475690
rect -960 475632 3330 475688
rect 3386 475632 3391 475688
rect -960 475630 3391 475632
rect -960 475540 480 475630
rect 3325 475627 3391 475630
rect 580533 471474 580599 471477
rect 583520 471474 584960 471564
rect 580533 471472 584960 471474
rect 580533 471416 580538 471472
rect 580594 471416 584960 471472
rect 580533 471414 584960 471416
rect 580533 471411 580599 471414
rect 583520 471324 584960 471414
rect -960 462634 480 462724
rect 3325 462634 3391 462637
rect -960 462632 3391 462634
rect -960 462576 3330 462632
rect 3386 462576 3391 462632
rect -960 462574 3391 462576
rect -960 462484 480 462574
rect 3325 462571 3391 462574
rect 579613 458146 579679 458149
rect 583520 458146 584960 458236
rect 579613 458144 584960 458146
rect 579613 458088 579618 458144
rect 579674 458088 584960 458144
rect 579613 458086 584960 458088
rect 579613 458083 579679 458086
rect 583520 457996 584960 458086
rect -960 449578 480 449668
rect 3325 449578 3391 449581
rect -960 449576 3391 449578
rect -960 449520 3330 449576
rect 3386 449520 3391 449576
rect -960 449518 3391 449520
rect -960 449428 480 449518
rect 3325 449515 3391 449518
rect 583520 444668 584960 444908
rect -960 436508 480 436748
rect 580441 431626 580507 431629
rect 583520 431626 584960 431716
rect 580441 431624 584960 431626
rect 580441 431568 580446 431624
rect 580502 431568 584960 431624
rect 580441 431566 584960 431568
rect 580441 431563 580507 431566
rect 583520 431476 584960 431566
rect -960 423602 480 423692
rect 3141 423602 3207 423605
rect -960 423600 3207 423602
rect -960 423544 3146 423600
rect 3202 423544 3207 423600
rect -960 423542 3207 423544
rect -960 423452 480 423542
rect 3141 423539 3207 423542
rect 579705 418298 579771 418301
rect 583520 418298 584960 418388
rect 579705 418296 584960 418298
rect 579705 418240 579710 418296
rect 579766 418240 584960 418296
rect 579705 418238 584960 418240
rect 579705 418235 579771 418238
rect 583520 418148 584960 418238
rect -960 410546 480 410636
rect 3693 410546 3759 410549
rect -960 410544 3759 410546
rect -960 410488 3698 410544
rect 3754 410488 3759 410544
rect -960 410486 3759 410488
rect -960 410396 480 410486
rect 3693 410483 3759 410486
rect 580165 404970 580231 404973
rect 583520 404970 584960 405060
rect 580165 404968 584960 404970
rect 580165 404912 580170 404968
rect 580226 404912 584960 404968
rect 580165 404910 584960 404912
rect 580165 404907 580231 404910
rect 583520 404820 584960 404910
rect -960 397490 480 397580
rect 3325 397490 3391 397493
rect -960 397488 3391 397490
rect -960 397432 3330 397488
rect 3386 397432 3391 397488
rect -960 397430 3391 397432
rect -960 397340 480 397430
rect 3325 397427 3391 397430
rect 583520 391628 584960 391868
rect -960 384284 480 384524
rect 580165 378450 580231 378453
rect 583520 378450 584960 378540
rect 580165 378448 584960 378450
rect 580165 378392 580170 378448
rect 580226 378392 584960 378448
rect 580165 378390 584960 378392
rect 580165 378387 580231 378390
rect 583520 378300 584960 378390
rect 38377 376954 38443 376957
rect 337653 376954 337719 376957
rect 38377 376952 39498 376954
rect 38377 376896 38382 376952
rect 38438 376924 39498 376952
rect 337653 376952 339418 376954
rect 38438 376896 40020 376924
rect 38377 376894 40020 376896
rect 38377 376891 38443 376894
rect 39438 376864 40020 376894
rect 337653 376896 337658 376952
rect 337714 376924 339418 376952
rect 337714 376896 340032 376924
rect 337653 376894 340032 376896
rect 337653 376891 337719 376894
rect 339358 376864 340032 376894
rect 37549 376002 37615 376005
rect 337745 376002 337811 376005
rect 37549 376000 39498 376002
rect 37549 375944 37554 376000
rect 37610 375972 39498 376000
rect 337745 376000 339418 376002
rect 37610 375944 40020 375972
rect 37549 375942 40020 375944
rect 37549 375939 37615 375942
rect 39438 375912 40020 375942
rect 337745 375944 337750 376000
rect 337806 375972 339418 376000
rect 337806 375944 340032 375972
rect 337745 375942 340032 375944
rect 337745 375939 337811 375942
rect 339358 375912 340032 375942
rect 38745 373826 38811 373829
rect 337469 373826 337535 373829
rect 38745 373824 39498 373826
rect 38745 373768 38750 373824
rect 38806 373796 39498 373824
rect 337469 373824 339418 373826
rect 38806 373768 40020 373796
rect 38745 373766 40020 373768
rect 38745 373763 38811 373766
rect 39438 373736 40020 373766
rect 337469 373768 337474 373824
rect 337530 373796 339418 373824
rect 337530 373768 340032 373796
rect 337469 373766 340032 373768
rect 337469 373763 337535 373766
rect 339358 373736 340032 373766
rect 38469 372874 38535 372877
rect 337561 372874 337627 372877
rect 38469 372872 39498 372874
rect 38469 372816 38474 372872
rect 38530 372844 39498 372872
rect 337561 372872 339418 372874
rect 38530 372816 40020 372844
rect 38469 372814 40020 372816
rect 38469 372811 38535 372814
rect 39438 372784 40020 372814
rect 337561 372816 337566 372872
rect 337622 372844 339418 372872
rect 337622 372816 340032 372844
rect 337561 372814 340032 372816
rect 337561 372811 337627 372814
rect 339358 372784 340032 372814
rect -960 371378 480 371468
rect 3325 371378 3391 371381
rect -960 371376 3391 371378
rect -960 371320 3330 371376
rect 3386 371320 3391 371376
rect -960 371318 3391 371320
rect -960 371228 480 371318
rect 3325 371315 3391 371318
rect 37917 371106 37983 371109
rect 337469 371106 337535 371109
rect 37917 371104 39498 371106
rect 37917 371048 37922 371104
rect 37978 371076 39498 371104
rect 337469 371104 339418 371106
rect 37978 371048 40020 371076
rect 37917 371046 40020 371048
rect 37917 371043 37983 371046
rect 39438 371016 40020 371046
rect 337469 371048 337474 371104
rect 337530 371076 339418 371104
rect 337530 371048 340032 371076
rect 337469 371046 340032 371048
rect 337469 371043 337535 371046
rect 339358 371016 340032 371046
rect 38653 370018 38719 370021
rect 337745 370018 337811 370021
rect 38653 370016 39498 370018
rect 38653 369960 38658 370016
rect 38714 369988 39498 370016
rect 337745 370016 339418 370018
rect 38714 369960 40020 369988
rect 38653 369958 40020 369960
rect 38653 369955 38719 369958
rect 39438 369928 40020 369958
rect 337745 369960 337750 370016
rect 337806 369988 339418 370016
rect 337806 369960 340032 369988
rect 337745 369958 340032 369960
rect 337745 369955 337811 369958
rect 339358 369928 340032 369958
rect 38837 368250 38903 368253
rect 337469 368250 337535 368253
rect 38837 368248 39498 368250
rect 38837 368192 38842 368248
rect 38898 368220 39498 368248
rect 337469 368248 339418 368250
rect 38898 368192 40020 368220
rect 38837 368190 40020 368192
rect 38837 368187 38903 368190
rect 39438 368160 40020 368190
rect 337469 368192 337474 368248
rect 337530 368220 339418 368248
rect 337530 368192 340032 368220
rect 337469 368190 340032 368192
rect 337469 368187 337535 368190
rect 339358 368160 340032 368190
rect 580165 365122 580231 365125
rect 583520 365122 584960 365212
rect 580165 365120 584960 365122
rect 580165 365064 580170 365120
rect 580226 365064 584960 365120
rect 580165 365062 584960 365064
rect 580165 365059 580231 365062
rect 583520 364972 584960 365062
rect -960 358458 480 358548
rect 3785 358458 3851 358461
rect -960 358456 3851 358458
rect -960 358400 3790 358456
rect 3846 358400 3851 358456
rect -960 358398 3851 358400
rect -960 358308 480 358398
rect 3785 358395 3851 358398
rect 580165 351930 580231 351933
rect 583520 351930 584960 352020
rect 580165 351928 584960 351930
rect 580165 351872 580170 351928
rect 580226 351872 584960 351928
rect 580165 351870 584960 351872
rect 580165 351867 580231 351870
rect 583520 351780 584960 351870
rect 38193 350026 38259 350029
rect 337745 350026 337811 350029
rect 38193 350024 39498 350026
rect 38193 349968 38198 350024
rect 38254 349996 39498 350024
rect 337745 350024 339418 350026
rect 38254 349968 40020 349996
rect 38193 349966 40020 349968
rect 38193 349963 38259 349966
rect 39438 349936 40020 349966
rect 337745 349968 337750 350024
rect 337806 349996 339418 350024
rect 337806 349968 340032 349996
rect 337745 349966 340032 349968
rect 337745 349963 337811 349966
rect 339358 349936 340032 349966
rect 38561 348394 38627 348397
rect 337377 348394 337443 348397
rect 38561 348392 39498 348394
rect 38561 348336 38566 348392
rect 38622 348364 39498 348392
rect 337377 348392 339418 348394
rect 38622 348336 40020 348364
rect 38561 348334 40020 348336
rect 38561 348331 38627 348334
rect 39438 348304 40020 348334
rect 337377 348336 337382 348392
rect 337438 348364 339418 348392
rect 337438 348336 340032 348364
rect 337377 348334 340032 348336
rect 337377 348331 337443 348334
rect 339358 348304 340032 348334
rect 37641 348122 37707 348125
rect 337653 348122 337719 348125
rect 37641 348120 39498 348122
rect 37641 348064 37646 348120
rect 37702 348092 39498 348120
rect 337653 348120 339418 348122
rect 37702 348064 40020 348092
rect 37641 348062 40020 348064
rect 37641 348059 37707 348062
rect 39438 348032 40020 348062
rect 337653 348064 337658 348120
rect 337714 348092 339418 348120
rect 337714 348064 340032 348092
rect 337653 348062 340032 348064
rect 337653 348059 337719 348062
rect 339358 348032 340032 348062
rect -960 345402 480 345492
rect 3049 345402 3115 345405
rect -960 345400 3115 345402
rect -960 345344 3054 345400
rect 3110 345344 3115 345400
rect -960 345342 3115 345344
rect -960 345252 480 345342
rect 3049 345339 3115 345342
rect 583520 338452 584960 338692
rect 76966 338132 76972 338196
rect 77036 338132 77042 338196
rect 80646 338132 80652 338196
rect 80716 338132 80722 338196
rect 83958 338132 83964 338196
rect 84028 338132 84034 338196
rect 90950 338132 90956 338196
rect 91020 338132 91026 338196
rect 98494 338132 98500 338196
rect 98564 338132 98570 338196
rect 131062 338132 131068 338196
rect 131132 338132 131138 338196
rect 372286 338132 372292 338196
rect 372356 338132 372362 338196
rect 382774 338132 382780 338196
rect 382844 338132 382850 338196
rect 386454 338132 386460 338196
rect 386524 338132 386530 338196
rect 408166 338132 408172 338196
rect 408236 338132 408242 338196
rect 57830 337996 57836 338060
rect 57900 338058 57906 338060
rect 70710 338058 70716 338060
rect 57900 337998 70716 338058
rect 57900 337996 57906 337998
rect 70710 337996 70716 337998
rect 70780 337996 70786 338060
rect 76974 338058 77034 338132
rect 77201 338058 77267 338061
rect 76974 338056 77267 338058
rect 76974 338000 77206 338056
rect 77262 338000 77267 338056
rect 76974 337998 77267 338000
rect 80654 338058 80714 338132
rect 83966 338061 84026 338132
rect 90958 338061 91018 338132
rect 81249 338058 81315 338061
rect 80654 338056 81315 338058
rect 80654 338000 81254 338056
rect 81310 338000 81315 338056
rect 80654 337998 81315 338000
rect 83966 338056 84075 338061
rect 83966 338000 84014 338056
rect 84070 338000 84075 338056
rect 83966 337998 84075 338000
rect 90958 338056 91067 338061
rect 90958 338000 91006 338056
rect 91062 338000 91067 338056
rect 90958 337998 91067 338000
rect 77201 337995 77267 337998
rect 81249 337995 81315 337998
rect 84009 337995 84075 337998
rect 91001 337995 91067 337998
rect 97993 338058 98059 338061
rect 98502 338058 98562 338132
rect 131070 338061 131130 338132
rect 97993 338056 98562 338058
rect 97993 338000 97998 338056
rect 98054 338000 98562 338056
rect 97993 337998 98562 338000
rect 131021 338056 131130 338061
rect 131021 338000 131026 338056
rect 131082 338000 131130 338056
rect 131021 337998 131130 338000
rect 371233 338058 371299 338061
rect 372294 338058 372354 338132
rect 371233 338056 372354 338058
rect 371233 338000 371238 338056
rect 371294 338000 372354 338056
rect 371233 337998 372354 338000
rect 382365 338058 382431 338061
rect 382782 338058 382842 338132
rect 386462 338061 386522 338132
rect 382365 338056 382842 338058
rect 382365 338000 382370 338056
rect 382426 338000 382842 338056
rect 382365 337998 382842 338000
rect 386413 338056 386522 338061
rect 386413 338000 386418 338056
rect 386474 338000 386522 338056
rect 386413 337998 386522 338000
rect 407113 338058 407179 338061
rect 408174 338058 408234 338132
rect 407113 338056 408234 338058
rect 407113 338000 407118 338056
rect 407174 338000 408234 338056
rect 407113 337998 408234 338000
rect 97993 337995 98059 337998
rect 131021 337995 131087 337998
rect 371233 337995 371299 337998
rect 382365 337995 382431 337998
rect 386413 337995 386479 337998
rect 407113 337995 407179 337998
rect 59353 337922 59419 337925
rect 60590 337922 60596 337924
rect 59353 337920 60596 337922
rect 59353 337864 59358 337920
rect 59414 337864 60596 337920
rect 59353 337862 60596 337864
rect 59353 337859 59419 337862
rect 60590 337860 60596 337862
rect 60660 337860 60666 337924
rect 73654 337922 73660 337924
rect 68142 337862 73660 337922
rect 55990 337724 55996 337788
rect 56060 337786 56066 337788
rect 56501 337786 56567 337789
rect 56060 337784 56567 337786
rect 56060 337728 56506 337784
rect 56562 337728 56567 337784
rect 56060 337726 56567 337728
rect 56060 337724 56066 337726
rect 56501 337723 56567 337726
rect 57094 337724 57100 337788
rect 57164 337786 57170 337788
rect 57881 337786 57947 337789
rect 57164 337784 57947 337786
rect 57164 337728 57886 337784
rect 57942 337728 57947 337784
rect 57164 337726 57947 337728
rect 57164 337724 57170 337726
rect 57881 337723 57947 337726
rect 59670 337724 59676 337788
rect 59740 337786 59746 337788
rect 60641 337786 60707 337789
rect 59740 337784 60707 337786
rect 59740 337728 60646 337784
rect 60702 337728 60707 337784
rect 59740 337726 60707 337728
rect 59740 337724 59746 337726
rect 60641 337723 60707 337726
rect 62113 337786 62179 337789
rect 63166 337786 63172 337788
rect 62113 337784 63172 337786
rect 62113 337728 62118 337784
rect 62174 337728 63172 337784
rect 62113 337726 63172 337728
rect 62113 337723 62179 337726
rect 63166 337724 63172 337726
rect 63236 337724 63242 337788
rect 64270 337724 64276 337788
rect 64340 337786 64346 337788
rect 64781 337786 64847 337789
rect 64340 337784 64847 337786
rect 64340 337728 64786 337784
rect 64842 337728 64847 337784
rect 64340 337726 64847 337728
rect 64340 337724 64346 337726
rect 64781 337723 64847 337726
rect 53598 337588 53604 337652
rect 53668 337650 53674 337652
rect 68142 337650 68202 337862
rect 73654 337860 73660 337862
rect 73724 337860 73730 337924
rect 78070 337860 78076 337924
rect 78140 337922 78146 337924
rect 78581 337922 78647 337925
rect 78140 337920 78647 337922
rect 78140 337864 78586 337920
rect 78642 337864 78647 337920
rect 78140 337862 78647 337864
rect 78140 337860 78146 337862
rect 78581 337859 78647 337862
rect 93342 337860 93348 337924
rect 93412 337922 93418 337924
rect 93577 337922 93643 337925
rect 93412 337920 93643 337922
rect 93412 337864 93582 337920
rect 93638 337864 93643 337920
rect 93412 337862 93643 337864
rect 93412 337860 93418 337862
rect 93577 337859 93643 337862
rect 375373 337922 375439 337925
rect 379513 337924 379579 337925
rect 376150 337922 376156 337924
rect 375373 337920 376156 337922
rect 375373 337864 375378 337920
rect 375434 337864 376156 337920
rect 375373 337862 376156 337864
rect 375373 337859 375439 337862
rect 376150 337860 376156 337862
rect 376220 337860 376226 337924
rect 379462 337860 379468 337924
rect 379532 337922 379579 337924
rect 394693 337922 394759 337925
rect 395654 337922 395660 337924
rect 379532 337920 379624 337922
rect 379574 337864 379624 337920
rect 379532 337862 379624 337864
rect 394693 337920 395660 337922
rect 394693 337864 394698 337920
rect 394754 337864 395660 337920
rect 394693 337862 395660 337864
rect 379532 337860 379579 337862
rect 379513 337859 379579 337860
rect 394693 337859 394759 337862
rect 395654 337860 395660 337862
rect 395724 337860 395730 337924
rect 397453 337922 397519 337925
rect 398046 337922 398052 337924
rect 397453 337920 398052 337922
rect 397453 337864 397458 337920
rect 397514 337864 398052 337920
rect 397453 337862 398052 337864
rect 397453 337859 397519 337862
rect 398046 337860 398052 337862
rect 398116 337860 398122 337924
rect 68318 337724 68324 337788
rect 68388 337786 68394 337788
rect 68829 337786 68895 337789
rect 68388 337784 68895 337786
rect 68388 337728 68834 337784
rect 68890 337728 68895 337784
rect 68388 337726 68895 337728
rect 68388 337724 68394 337726
rect 68829 337723 68895 337726
rect 69657 337786 69723 337789
rect 78438 337786 78444 337788
rect 69657 337784 78444 337786
rect 69657 337728 69662 337784
rect 69718 337728 78444 337784
rect 69657 337726 78444 337728
rect 69657 337723 69723 337726
rect 78438 337724 78444 337726
rect 78508 337724 78514 337788
rect 85982 337724 85988 337788
rect 86052 337786 86058 337788
rect 86861 337786 86927 337789
rect 86052 337784 86927 337786
rect 86052 337728 86866 337784
rect 86922 337728 86927 337784
rect 86052 337726 86927 337728
rect 86052 337724 86058 337726
rect 86861 337723 86927 337726
rect 87137 337786 87203 337789
rect 88190 337786 88196 337788
rect 87137 337784 88196 337786
rect 87137 337728 87142 337784
rect 87198 337728 88196 337784
rect 87137 337726 88196 337728
rect 87137 337723 87203 337726
rect 88190 337724 88196 337726
rect 88260 337724 88266 337788
rect 88742 337724 88748 337788
rect 88812 337786 88818 337788
rect 89621 337786 89687 337789
rect 88812 337784 89687 337786
rect 88812 337728 89626 337784
rect 89682 337728 89687 337784
rect 88812 337726 89687 337728
rect 88812 337724 88818 337726
rect 89621 337723 89687 337726
rect 91502 337724 91508 337788
rect 91572 337786 91578 337788
rect 92381 337786 92447 337789
rect 91572 337784 92447 337786
rect 91572 337728 92386 337784
rect 92442 337728 92447 337784
rect 91572 337726 92447 337728
rect 91572 337724 91578 337726
rect 92381 337723 92447 337726
rect 96613 337786 96679 337789
rect 97022 337786 97028 337788
rect 96613 337784 97028 337786
rect 96613 337728 96618 337784
rect 96674 337728 97028 337784
rect 96613 337726 97028 337728
rect 96613 337723 96679 337726
rect 97022 337724 97028 337726
rect 97092 337724 97098 337788
rect 103278 337724 103284 337788
rect 103348 337786 103354 337788
rect 104801 337786 104867 337789
rect 103348 337784 104867 337786
rect 103348 337728 104806 337784
rect 104862 337728 104867 337784
rect 103348 337726 104867 337728
rect 103348 337724 103354 337726
rect 104801 337723 104867 337726
rect 113173 337786 113239 337789
rect 113398 337786 113404 337788
rect 113173 337784 113404 337786
rect 113173 337728 113178 337784
rect 113234 337728 113404 337784
rect 113173 337726 113404 337728
rect 113173 337723 113239 337726
rect 113398 337724 113404 337726
rect 113468 337724 113474 337788
rect 115974 337724 115980 337788
rect 116044 337786 116050 337788
rect 117221 337786 117287 337789
rect 118601 337788 118667 337789
rect 116044 337784 117287 337786
rect 116044 337728 117226 337784
rect 117282 337728 117287 337784
rect 116044 337726 117287 337728
rect 116044 337724 116050 337726
rect 117221 337723 117287 337726
rect 118550 337724 118556 337788
rect 118620 337786 118667 337788
rect 122833 337786 122899 337789
rect 123518 337786 123524 337788
rect 118620 337784 118712 337786
rect 118662 337728 118712 337784
rect 118620 337726 118712 337728
rect 122833 337784 123524 337786
rect 122833 337728 122838 337784
rect 122894 337728 123524 337784
rect 122833 337726 123524 337728
rect 118620 337724 118667 337726
rect 118601 337723 118667 337724
rect 122833 337723 122899 337726
rect 123518 337724 123524 337726
rect 123588 337724 123594 337788
rect 125593 337786 125659 337789
rect 125910 337786 125916 337788
rect 125593 337784 125916 337786
rect 125593 337728 125598 337784
rect 125654 337728 125916 337784
rect 125593 337726 125916 337728
rect 125593 337723 125659 337726
rect 125910 337724 125916 337726
rect 125980 337724 125986 337788
rect 133454 337724 133460 337788
rect 133524 337786 133530 337788
rect 133781 337786 133847 337789
rect 133524 337784 133847 337786
rect 133524 337728 133786 337784
rect 133842 337728 133847 337784
rect 133524 337726 133847 337728
rect 133524 337724 133530 337726
rect 133781 337723 133847 337726
rect 135846 337724 135852 337788
rect 135916 337786 135922 337788
rect 136541 337786 136607 337789
rect 135916 337784 136607 337786
rect 135916 337728 136546 337784
rect 136602 337728 136607 337784
rect 135916 337726 136607 337728
rect 135916 337724 135922 337726
rect 136541 337723 136607 337726
rect 138606 337724 138612 337788
rect 138676 337786 138682 337788
rect 139301 337786 139367 337789
rect 143441 337788 143507 337789
rect 138676 337784 139367 337786
rect 138676 337728 139306 337784
rect 139362 337728 139367 337784
rect 138676 337726 139367 337728
rect 138676 337724 138682 337726
rect 139301 337723 139367 337726
rect 143390 337724 143396 337788
rect 143460 337786 143507 337788
rect 143460 337784 143552 337786
rect 143502 337728 143552 337784
rect 143460 337726 143552 337728
rect 143460 337724 143507 337726
rect 145966 337724 145972 337788
rect 146036 337786 146042 337788
rect 146201 337786 146267 337789
rect 146036 337784 146267 337786
rect 146036 337728 146206 337784
rect 146262 337728 146267 337784
rect 146036 337726 146267 337728
rect 146036 337724 146042 337726
rect 143441 337723 143507 337724
rect 146201 337723 146267 337726
rect 362953 337786 363019 337789
rect 364190 337786 364196 337788
rect 362953 337784 364196 337786
rect 362953 337728 362958 337784
rect 363014 337728 364196 337784
rect 362953 337726 364196 337728
rect 362953 337723 363019 337726
rect 364190 337724 364196 337726
rect 364260 337724 364266 337788
rect 366357 337786 366423 337789
rect 367502 337786 367508 337788
rect 366357 337784 367508 337786
rect 366357 337728 366362 337784
rect 366418 337728 367508 337784
rect 366357 337726 367508 337728
rect 366357 337723 366423 337726
rect 367502 337724 367508 337726
rect 367572 337724 367578 337788
rect 369853 337786 369919 337789
rect 370078 337786 370084 337788
rect 369853 337784 370084 337786
rect 369853 337728 369858 337784
rect 369914 337728 370084 337784
rect 369853 337726 370084 337728
rect 369853 337723 369919 337726
rect 370078 337724 370084 337726
rect 370148 337724 370154 337788
rect 372613 337786 372679 337789
rect 373574 337786 373580 337788
rect 372613 337784 373580 337786
rect 372613 337728 372618 337784
rect 372674 337728 373580 337784
rect 372613 337726 373580 337728
rect 372613 337723 372679 337726
rect 373574 337724 373580 337726
rect 373644 337724 373650 337788
rect 378133 337786 378199 337789
rect 378542 337786 378548 337788
rect 378133 337784 378548 337786
rect 378133 337728 378138 337784
rect 378194 337728 378548 337784
rect 378133 337726 378548 337728
rect 378133 337723 378199 337726
rect 378542 337724 378548 337726
rect 378612 337724 378618 337788
rect 380157 337786 380223 337789
rect 381670 337786 381676 337788
rect 380157 337784 381676 337786
rect 380157 337728 380162 337784
rect 380218 337728 381676 337784
rect 380157 337726 381676 337728
rect 380157 337723 380223 337726
rect 381670 337724 381676 337726
rect 381740 337724 381746 337788
rect 389173 337786 389239 337789
rect 389766 337786 389772 337788
rect 389173 337784 389772 337786
rect 389173 337728 389178 337784
rect 389234 337728 389772 337784
rect 389173 337726 389772 337728
rect 389173 337723 389239 337726
rect 389766 337724 389772 337726
rect 389836 337724 389842 337788
rect 391933 337786 391999 337789
rect 392158 337786 392164 337788
rect 391933 337784 392164 337786
rect 391933 337728 391938 337784
rect 391994 337728 392164 337784
rect 391933 337726 392164 337728
rect 391933 337723 391999 337726
rect 392158 337724 392164 337726
rect 392228 337724 392234 337788
rect 53668 337590 68202 337650
rect 53668 337588 53674 337590
rect 68686 337588 68692 337652
rect 68756 337650 68762 337652
rect 68921 337650 68987 337653
rect 71313 337652 71379 337653
rect 74625 337652 74691 337653
rect 68756 337648 68987 337650
rect 68756 337592 68926 337648
rect 68982 337592 68987 337648
rect 68756 337590 68987 337592
rect 68756 337588 68762 337590
rect 68921 337587 68987 337590
rect 71262 337588 71268 337652
rect 71332 337650 71379 337652
rect 71332 337648 71424 337650
rect 71374 337592 71424 337648
rect 71332 337590 71424 337592
rect 71332 337588 71379 337590
rect 74574 337588 74580 337652
rect 74644 337650 74691 337652
rect 74644 337648 74736 337650
rect 74686 337592 74736 337648
rect 74644 337590 74736 337592
rect 74644 337588 74691 337590
rect 79542 337588 79548 337652
rect 79612 337650 79618 337652
rect 79961 337650 80027 337653
rect 79612 337648 80027 337650
rect 79612 337592 79966 337648
rect 80022 337592 80027 337648
rect 79612 337590 80027 337592
rect 79612 337588 79618 337590
rect 71313 337587 71379 337588
rect 74625 337587 74691 337588
rect 79961 337587 80027 337590
rect 81750 337588 81756 337652
rect 81820 337650 81826 337652
rect 82169 337650 82235 337653
rect 81820 337648 82235 337650
rect 81820 337592 82174 337648
rect 82230 337592 82235 337648
rect 81820 337590 82235 337592
rect 81820 337588 81826 337590
rect 82169 337587 82235 337590
rect 82905 337650 82971 337653
rect 83406 337650 83412 337652
rect 82905 337648 83412 337650
rect 82905 337592 82910 337648
rect 82966 337592 83412 337648
rect 82905 337590 83412 337592
rect 82905 337587 82971 337590
rect 83406 337588 83412 337590
rect 83476 337588 83482 337652
rect 85246 337588 85252 337652
rect 85316 337650 85322 337652
rect 85481 337650 85547 337653
rect 85316 337648 85547 337650
rect 85316 337592 85486 337648
rect 85542 337592 85547 337648
rect 85316 337590 85547 337592
rect 85316 337588 85322 337590
rect 85481 337587 85547 337590
rect 85665 337650 85731 337653
rect 86350 337650 86356 337652
rect 85665 337648 86356 337650
rect 85665 337592 85670 337648
rect 85726 337592 86356 337648
rect 85665 337590 86356 337592
rect 85665 337587 85731 337590
rect 86350 337588 86356 337590
rect 86420 337588 86426 337652
rect 87045 337650 87111 337653
rect 87638 337650 87644 337652
rect 87045 337648 87644 337650
rect 87045 337592 87050 337648
rect 87106 337592 87644 337648
rect 87045 337590 87644 337592
rect 87045 337587 87111 337590
rect 87638 337588 87644 337590
rect 87708 337588 87714 337652
rect 89713 337650 89779 337653
rect 89846 337650 89852 337652
rect 89713 337648 89852 337650
rect 89713 337592 89718 337648
rect 89774 337592 89852 337648
rect 89713 337590 89852 337592
rect 89713 337587 89779 337590
rect 89846 337588 89852 337590
rect 89916 337588 89922 337652
rect 91185 337650 91251 337653
rect 92238 337650 92244 337652
rect 91185 337648 92244 337650
rect 91185 337592 91190 337648
rect 91246 337592 92244 337648
rect 91185 337590 92244 337592
rect 91185 337587 91251 337590
rect 92238 337588 92244 337590
rect 92308 337588 92314 337652
rect 93526 337588 93532 337652
rect 93596 337650 93602 337652
rect 93669 337650 93735 337653
rect 93596 337648 93735 337650
rect 93596 337592 93674 337648
rect 93730 337592 93735 337648
rect 93596 337590 93735 337592
rect 93596 337588 93602 337590
rect 93669 337587 93735 337590
rect 95734 337588 95740 337652
rect 95804 337650 95810 337652
rect 96337 337650 96403 337653
rect 95804 337648 96403 337650
rect 95804 337592 96342 337648
rect 96398 337592 96403 337648
rect 95804 337590 96403 337592
rect 95804 337588 95810 337590
rect 96337 337587 96403 337590
rect 97942 337588 97948 337652
rect 98012 337650 98018 337652
rect 99097 337650 99163 337653
rect 99281 337652 99347 337653
rect 98012 337648 99163 337650
rect 98012 337592 99102 337648
rect 99158 337592 99163 337648
rect 98012 337590 99163 337592
rect 98012 337588 98018 337590
rect 99097 337587 99163 337590
rect 99230 337588 99236 337652
rect 99300 337650 99347 337652
rect 99300 337648 99392 337650
rect 99342 337592 99392 337648
rect 99300 337590 99392 337592
rect 99300 337588 99347 337590
rect 100886 337588 100892 337652
rect 100956 337650 100962 337652
rect 102041 337650 102107 337653
rect 100956 337648 102107 337650
rect 100956 337592 102046 337648
rect 102102 337592 102107 337648
rect 100956 337590 102107 337592
rect 100956 337588 100962 337590
rect 99281 337587 99347 337588
rect 102041 337587 102107 337590
rect 104893 337650 104959 337653
rect 105854 337650 105860 337652
rect 104893 337648 105860 337650
rect 104893 337592 104898 337648
rect 104954 337592 105860 337648
rect 104893 337590 105860 337592
rect 104893 337587 104959 337590
rect 105854 337588 105860 337590
rect 105924 337588 105930 337652
rect 108246 337588 108252 337652
rect 108316 337650 108322 337652
rect 108941 337650 109007 337653
rect 108316 337648 109007 337650
rect 108316 337592 108946 337648
rect 109002 337592 109007 337648
rect 108316 337590 109007 337592
rect 108316 337588 108322 337590
rect 108941 337587 109007 337590
rect 111006 337588 111012 337652
rect 111076 337650 111082 337652
rect 233182 337650 233188 337652
rect 111076 337590 233188 337650
rect 111076 337588 111082 337590
rect 233182 337588 233188 337590
rect 233252 337588 233258 337652
rect 356053 337650 356119 337653
rect 357014 337650 357020 337652
rect 356053 337648 357020 337650
rect 356053 337592 356058 337648
rect 356114 337592 357020 337648
rect 356053 337590 357020 337592
rect 356053 337587 356119 337590
rect 357014 337588 357020 337590
rect 357084 337588 357090 337652
rect 357433 337650 357499 337653
rect 358118 337650 358124 337652
rect 357433 337648 358124 337650
rect 357433 337592 357438 337648
rect 357494 337592 358124 337648
rect 357433 337590 358124 337592
rect 357433 337587 357499 337590
rect 358118 337588 358124 337590
rect 358188 337588 358194 337652
rect 358813 337650 358879 337653
rect 359590 337650 359596 337652
rect 358813 337648 359596 337650
rect 358813 337592 358818 337648
rect 358874 337592 359596 337648
rect 358813 337590 359596 337592
rect 358813 337587 358879 337590
rect 359590 337588 359596 337590
rect 359660 337588 359666 337652
rect 360193 337650 360259 337653
rect 360510 337650 360516 337652
rect 360193 337648 360516 337650
rect 360193 337592 360198 337648
rect 360254 337592 360516 337648
rect 360193 337590 360516 337592
rect 360193 337587 360259 337590
rect 360510 337588 360516 337590
rect 360580 337588 360586 337652
rect 361573 337650 361639 337653
rect 363045 337652 363111 337653
rect 361798 337650 361804 337652
rect 361573 337648 361804 337650
rect 361573 337592 361578 337648
rect 361634 337592 361804 337648
rect 361573 337590 361804 337592
rect 361573 337587 361639 337590
rect 361798 337588 361804 337590
rect 361868 337588 361874 337652
rect 363045 337650 363092 337652
rect 363000 337648 363092 337650
rect 363000 337592 363050 337648
rect 363000 337590 363092 337592
rect 363045 337588 363092 337590
rect 363156 337588 363162 337652
rect 365713 337650 365779 337653
rect 366398 337650 366404 337652
rect 365713 337648 366404 337650
rect 365713 337592 365718 337648
rect 365774 337592 366404 337648
rect 365713 337590 366404 337592
rect 363045 337587 363111 337588
rect 365713 337587 365779 337590
rect 366398 337588 366404 337590
rect 366468 337588 366474 337652
rect 367185 337650 367251 337653
rect 368054 337650 368060 337652
rect 367185 337648 368060 337650
rect 367185 337592 367190 337648
rect 367246 337592 368060 337648
rect 367185 337590 368060 337592
rect 367185 337587 367251 337590
rect 368054 337588 368060 337590
rect 368124 337588 368130 337652
rect 368473 337650 368539 337653
rect 368974 337650 368980 337652
rect 368473 337648 368980 337650
rect 368473 337592 368478 337648
rect 368534 337592 368980 337648
rect 368473 337590 368980 337592
rect 368473 337587 368539 337590
rect 368974 337588 368980 337590
rect 369044 337588 369050 337652
rect 369945 337650 370011 337653
rect 370630 337650 370636 337652
rect 369945 337648 370636 337650
rect 369945 337592 369950 337648
rect 370006 337592 370636 337648
rect 369945 337590 370636 337592
rect 369945 337587 370011 337590
rect 370630 337588 370636 337590
rect 370700 337588 370706 337652
rect 371877 337650 371943 337653
rect 373390 337650 373396 337652
rect 371877 337648 373396 337650
rect 371877 337592 371882 337648
rect 371938 337592 373396 337648
rect 371877 337590 373396 337592
rect 371877 337587 371943 337590
rect 373390 337588 373396 337590
rect 373460 337588 373466 337652
rect 373993 337650 374059 337653
rect 374494 337650 374500 337652
rect 373993 337648 374500 337650
rect 373993 337592 373998 337648
rect 374054 337592 374500 337648
rect 373993 337590 374500 337592
rect 373993 337587 374059 337590
rect 374494 337588 374500 337590
rect 374564 337588 374570 337652
rect 375465 337650 375531 337653
rect 375782 337650 375788 337652
rect 375465 337648 375788 337650
rect 375465 337592 375470 337648
rect 375526 337592 375788 337648
rect 375465 337590 375788 337592
rect 375465 337587 375531 337590
rect 375782 337588 375788 337590
rect 375852 337588 375858 337652
rect 376753 337650 376819 337653
rect 377990 337650 377996 337652
rect 376753 337648 377996 337650
rect 376753 337592 376758 337648
rect 376814 337592 377996 337648
rect 376753 337590 377996 337592
rect 376753 337587 376819 337590
rect 377990 337588 377996 337590
rect 378060 337588 378066 337652
rect 380985 337650 381051 337653
rect 381118 337650 381124 337652
rect 380985 337648 381124 337650
rect 380985 337592 380990 337648
rect 381046 337592 381124 337648
rect 380985 337590 381124 337592
rect 380985 337587 381051 337590
rect 381118 337588 381124 337590
rect 381188 337588 381194 337652
rect 384297 337650 384363 337653
rect 385166 337650 385172 337652
rect 384297 337648 385172 337650
rect 384297 337592 384302 337648
rect 384358 337592 385172 337648
rect 384297 337590 385172 337592
rect 384297 337587 384363 337590
rect 385166 337588 385172 337590
rect 385236 337588 385242 337652
rect 390553 337650 390619 337653
rect 393405 337652 393471 337653
rect 391054 337650 391060 337652
rect 390553 337648 391060 337650
rect 390553 337592 390558 337648
rect 390614 337592 391060 337648
rect 390553 337590 391060 337592
rect 390553 337587 390619 337590
rect 391054 337588 391060 337590
rect 391124 337588 391130 337652
rect 393405 337650 393452 337652
rect 393360 337648 393452 337650
rect 393360 337592 393410 337648
rect 393360 337590 393452 337592
rect 393405 337588 393452 337590
rect 393516 337588 393522 337652
rect 395337 337650 395403 337653
rect 396022 337650 396028 337652
rect 395337 337648 396028 337650
rect 395337 337592 395342 337648
rect 395398 337592 396028 337648
rect 395337 337590 396028 337592
rect 393405 337587 393471 337588
rect 395337 337587 395403 337590
rect 396022 337588 396028 337590
rect 396092 337588 396098 337652
rect 398097 337650 398163 337653
rect 399150 337650 399156 337652
rect 398097 337648 399156 337650
rect 398097 337592 398102 337648
rect 398158 337592 399156 337648
rect 398097 337590 399156 337592
rect 398097 337587 398163 337590
rect 399150 337588 399156 337590
rect 399220 337588 399226 337652
rect 399569 337650 399635 337653
rect 401174 337650 401180 337652
rect 399569 337648 401180 337650
rect 399569 337592 399574 337648
rect 399630 337592 401180 337648
rect 399569 337590 401180 337592
rect 399569 337587 399635 337590
rect 401174 337588 401180 337590
rect 401244 337588 401250 337652
rect 412633 337650 412699 337653
rect 413318 337650 413324 337652
rect 412633 337648 413324 337650
rect 412633 337592 412638 337648
rect 412694 337592 413324 337648
rect 412633 337590 413324 337592
rect 412633 337587 412699 337590
rect 413318 337588 413324 337590
rect 413388 337588 413394 337652
rect 415393 337650 415459 337653
rect 415894 337650 415900 337652
rect 415393 337648 415900 337650
rect 415393 337592 415398 337648
rect 415454 337592 415900 337648
rect 415393 337590 415900 337592
rect 415393 337587 415459 337590
rect 415894 337588 415900 337590
rect 415964 337588 415970 337652
rect 417417 337650 417483 337653
rect 420913 337652 420979 337653
rect 418286 337650 418292 337652
rect 417417 337648 418292 337650
rect 417417 337592 417422 337648
rect 417478 337592 418292 337648
rect 417417 337590 418292 337592
rect 417417 337587 417483 337590
rect 418286 337588 418292 337590
rect 418356 337588 418362 337652
rect 420862 337588 420868 337652
rect 420932 337650 420979 337652
rect 427813 337650 427879 337653
rect 428590 337650 428596 337652
rect 420932 337648 421024 337650
rect 420974 337592 421024 337648
rect 420932 337590 421024 337592
rect 427813 337648 428596 337650
rect 427813 337592 427818 337648
rect 427874 337592 428596 337648
rect 427813 337590 428596 337592
rect 420932 337588 420979 337590
rect 420913 337587 420979 337588
rect 427813 337587 427879 337590
rect 428590 337588 428596 337590
rect 428660 337588 428666 337652
rect 430573 337650 430639 337653
rect 430982 337650 430988 337652
rect 430573 337648 430988 337650
rect 430573 337592 430578 337648
rect 430634 337592 430988 337648
rect 430573 337590 430988 337592
rect 430573 337587 430639 337590
rect 430982 337588 430988 337590
rect 431052 337588 431058 337652
rect 434713 337650 434779 337653
rect 435766 337650 435772 337652
rect 434713 337648 435772 337650
rect 434713 337592 434718 337648
rect 434774 337592 435772 337648
rect 434713 337590 435772 337592
rect 434713 337587 434779 337590
rect 435766 337588 435772 337590
rect 435836 337588 435842 337652
rect 437473 337650 437539 337653
rect 438342 337650 438348 337652
rect 437473 337648 438348 337650
rect 437473 337592 437478 337648
rect 437534 337592 438348 337648
rect 437473 337590 438348 337592
rect 437473 337587 437539 337590
rect 438342 337588 438348 337590
rect 438412 337588 438418 337652
rect 445753 337650 445819 337653
rect 445886 337650 445892 337652
rect 445753 337648 445892 337650
rect 445753 337592 445758 337648
rect 445814 337592 445892 337648
rect 445753 337590 445892 337592
rect 445753 337587 445819 337590
rect 445886 337588 445892 337590
rect 445956 337588 445962 337652
rect 57973 337514 58039 337517
rect 58198 337514 58204 337516
rect 57973 337512 58204 337514
rect 57973 337456 57978 337512
rect 58034 337456 58204 337512
rect 57973 337454 58204 337456
rect 57973 337451 58039 337454
rect 58198 337452 58204 337454
rect 58268 337452 58274 337516
rect 59997 337514 60063 337517
rect 72366 337514 72372 337516
rect 59997 337512 72372 337514
rect 59997 337456 60002 337512
rect 60058 337456 72372 337512
rect 59997 337454 72372 337456
rect 59997 337451 60063 337454
rect 72366 337452 72372 337454
rect 72436 337452 72442 337516
rect 81014 337452 81020 337516
rect 81084 337514 81090 337516
rect 81341 337514 81407 337517
rect 81084 337512 81407 337514
rect 81084 337456 81346 337512
rect 81402 337456 81407 337512
rect 81084 337454 81407 337456
rect 81084 337452 81090 337454
rect 81341 337451 81407 337454
rect 82854 337452 82860 337516
rect 82924 337514 82930 337516
rect 231894 337514 231900 337516
rect 82924 337454 231900 337514
rect 82924 337452 82930 337454
rect 231894 337452 231900 337454
rect 231964 337452 231970 337516
rect 385033 337514 385099 337517
rect 385902 337514 385908 337516
rect 385033 337512 385908 337514
rect 385033 337456 385038 337512
rect 385094 337456 385908 337512
rect 385033 337454 385908 337456
rect 385033 337451 385099 337454
rect 385902 337452 385908 337454
rect 385972 337452 385978 337516
rect 387793 337514 387859 337517
rect 388294 337514 388300 337516
rect 387793 337512 388300 337514
rect 387793 337456 387798 337512
rect 387854 337456 388300 337512
rect 387793 337454 388300 337456
rect 387793 337451 387859 337454
rect 388294 337452 388300 337454
rect 388364 337452 388370 337516
rect 40401 337378 40467 337381
rect 356094 337378 356100 337380
rect 40401 337376 356100 337378
rect 40401 337320 40406 337376
rect 40462 337320 356100 337376
rect 40401 337318 356100 337320
rect 40401 337315 40467 337318
rect 356094 337316 356100 337318
rect 356164 337316 356170 337380
rect 382273 337378 382339 337381
rect 383510 337378 383516 337380
rect 382273 337376 383516 337378
rect 382273 337320 382278 337376
rect 382334 337320 383516 337376
rect 382273 337318 383516 337320
rect 382273 337315 382339 337318
rect 383510 337316 383516 337318
rect 383580 337316 383586 337380
rect 422937 337378 423003 337381
rect 423438 337378 423444 337380
rect 422937 337376 423444 337378
rect 422937 337320 422942 337376
rect 422998 337320 423444 337376
rect 422937 337318 423444 337320
rect 422937 337315 423003 337318
rect 423438 337316 423444 337318
rect 423508 337316 423514 337380
rect 52310 337180 52316 337244
rect 52380 337242 52386 337244
rect 59997 337242 60063 337245
rect 52380 337240 60063 337242
rect 52380 337184 60002 337240
rect 60058 337184 60063 337240
rect 52380 337182 60063 337184
rect 52380 337180 52386 337182
rect 59997 337179 60063 337182
rect 60733 337242 60799 337245
rect 61694 337242 61700 337244
rect 60733 337240 61700 337242
rect 60733 337184 60738 337240
rect 60794 337184 61700 337240
rect 60733 337182 61700 337184
rect 60733 337179 60799 337182
rect 61694 337180 61700 337182
rect 61764 337180 61770 337244
rect 65374 337180 65380 337244
rect 65444 337242 65450 337244
rect 66161 337242 66227 337245
rect 65444 337240 66227 337242
rect 65444 337184 66166 337240
rect 66222 337184 66227 337240
rect 65444 337182 66227 337184
rect 65444 337180 65450 337182
rect 66161 337179 66227 337182
rect 66662 337180 66668 337244
rect 66732 337242 66738 337244
rect 67541 337242 67607 337245
rect 66732 337240 67607 337242
rect 66732 337184 67546 337240
rect 67602 337184 67607 337240
rect 66732 337182 67607 337184
rect 66732 337180 66738 337182
rect 67541 337179 67607 337182
rect 386505 337242 386571 337245
rect 387558 337242 387564 337244
rect 386505 337240 387564 337242
rect 386505 337184 386510 337240
rect 386566 337184 387564 337240
rect 386505 337182 387564 337184
rect 386505 337179 386571 337182
rect 387558 337180 387564 337182
rect 387628 337180 387634 337244
rect 409873 337242 409939 337245
rect 410926 337242 410932 337244
rect 409873 337240 410932 337242
rect 409873 337184 409878 337240
rect 409934 337184 410932 337240
rect 409873 337182 410932 337184
rect 409873 337179 409939 337182
rect 410926 337180 410932 337182
rect 410996 337180 411002 337244
rect 442993 337242 443059 337245
rect 443310 337242 443316 337244
rect 442993 337240 443316 337242
rect 442993 337184 442998 337240
rect 443054 337184 443316 337240
rect 442993 337182 443316 337184
rect 442993 337179 443059 337182
rect 443310 337180 443316 337182
rect 443380 337180 443386 337244
rect 56358 337044 56364 337108
rect 56428 337106 56434 337108
rect 67582 337106 67588 337108
rect 56428 337046 67588 337106
rect 56428 337044 56434 337046
rect 67582 337044 67588 337046
rect 67652 337044 67658 337108
rect 140998 337044 141004 337108
rect 141068 337106 141074 337108
rect 142061 337106 142127 337109
rect 141068 337104 142127 337106
rect 141068 337048 142066 337104
rect 142122 337048 142127 337104
rect 141068 337046 142127 337048
rect 141068 337044 141074 337046
rect 142061 337043 142127 337046
rect 379513 337106 379579 337109
rect 380566 337106 380572 337108
rect 379513 337104 380572 337106
rect 379513 337048 379518 337104
rect 379574 337048 380572 337104
rect 379513 337046 380572 337048
rect 379513 337043 379579 337046
rect 380566 337044 380572 337046
rect 380636 337044 380642 337108
rect 387793 337106 387859 337109
rect 388662 337106 388668 337108
rect 387793 337104 388668 337106
rect 387793 337048 387798 337104
rect 387854 337048 388668 337104
rect 387793 337046 388668 337048
rect 387793 337043 387859 337046
rect 388662 337044 388668 337046
rect 388732 337044 388738 337108
rect 392577 337106 392643 337109
rect 394366 337106 394372 337108
rect 392577 337104 394372 337106
rect 392577 337048 392582 337104
rect 392638 337048 394372 337104
rect 392577 337046 394372 337048
rect 392577 337043 392643 337046
rect 394366 337044 394372 337046
rect 394436 337044 394442 337108
rect 433333 337106 433399 337109
rect 433558 337106 433564 337108
rect 433333 337104 433564 337106
rect 433333 337048 433338 337104
rect 433394 337048 433564 337104
rect 433333 337046 433564 337048
rect 433333 337043 433399 337046
rect 433558 337044 433564 337046
rect 433628 337044 433634 337108
rect 440233 337106 440299 337109
rect 440918 337106 440924 337108
rect 440233 337104 440924 337106
rect 440233 337048 440238 337104
rect 440294 337048 440924 337104
rect 440233 337046 440924 337048
rect 440233 337043 440299 337046
rect 440918 337044 440924 337046
rect 440988 337044 440994 337108
rect 58198 336908 58204 336972
rect 58268 336970 58274 336972
rect 69657 336970 69723 336973
rect 58268 336968 69723 336970
rect 58268 336912 69662 336968
rect 69718 336912 69723 336968
rect 58268 336910 69723 336912
rect 58268 336908 58274 336910
rect 69657 336907 69723 336910
rect 383745 336970 383811 336973
rect 383878 336970 383884 336972
rect 383745 336968 383884 336970
rect 383745 336912 383750 336968
rect 383806 336912 383884 336968
rect 383745 336910 383884 336912
rect 383745 336907 383811 336910
rect 383878 336908 383884 336910
rect 383948 336908 383954 336972
rect 393078 336908 393084 336972
rect 393148 336970 393154 336972
rect 393313 336970 393379 336973
rect 393148 336968 393379 336970
rect 393148 336912 393318 336968
rect 393374 336912 393379 336968
rect 393148 336910 393379 336912
rect 393148 336908 393154 336910
rect 393313 336907 393379 336910
rect 396073 336970 396139 336973
rect 396574 336970 396580 336972
rect 396073 336968 396580 336970
rect 396073 336912 396078 336968
rect 396134 336912 396580 336968
rect 396073 336910 396580 336912
rect 396073 336907 396139 336910
rect 396574 336908 396580 336910
rect 396644 336908 396650 336972
rect 405733 336970 405799 336973
rect 405958 336970 405964 336972
rect 405733 336968 405964 336970
rect 405733 336912 405738 336968
rect 405794 336912 405964 336968
rect 405733 336910 405964 336912
rect 405733 336907 405799 336910
rect 405958 336908 405964 336910
rect 406028 336908 406034 336972
rect 425053 336970 425119 336973
rect 425646 336970 425652 336972
rect 425053 336968 425652 336970
rect 425053 336912 425058 336968
rect 425114 336912 425652 336968
rect 425053 336910 425652 336912
rect 425053 336907 425119 336910
rect 425646 336908 425652 336910
rect 425716 336908 425722 336972
rect 70158 336772 70164 336836
rect 70228 336834 70234 336836
rect 70301 336834 70367 336837
rect 70228 336832 70367 336834
rect 70228 336776 70306 336832
rect 70362 336776 70367 336832
rect 70228 336774 70367 336776
rect 70228 336772 70234 336774
rect 70301 336771 70367 336774
rect 75913 336834 75979 336837
rect 76046 336834 76052 336836
rect 75913 336832 76052 336834
rect 75913 336776 75918 336832
rect 75974 336776 76052 336832
rect 75913 336774 76052 336776
rect 75913 336771 75979 336774
rect 76046 336772 76052 336774
rect 76116 336772 76122 336836
rect 94262 336772 94268 336836
rect 94332 336834 94338 336836
rect 95141 336834 95207 336837
rect 94332 336832 95207 336834
rect 94332 336776 95146 336832
rect 95202 336776 95207 336832
rect 94332 336774 95207 336776
rect 94332 336772 94338 336774
rect 95141 336771 95207 336774
rect 96102 336772 96108 336836
rect 96172 336834 96178 336836
rect 96521 336834 96587 336837
rect 96172 336832 96587 336834
rect 96172 336776 96526 336832
rect 96582 336776 96587 336832
rect 96172 336774 96587 336776
rect 96172 336772 96178 336774
rect 96521 336771 96587 336774
rect 120942 336772 120948 336836
rect 121012 336834 121018 336836
rect 121269 336834 121335 336837
rect 121012 336832 121335 336834
rect 121012 336776 121274 336832
rect 121330 336776 121335 336832
rect 121012 336774 121335 336776
rect 121012 336772 121018 336774
rect 121269 336771 121335 336774
rect 128486 336772 128492 336836
rect 128556 336834 128562 336836
rect 129641 336834 129707 336837
rect 128556 336832 129707 336834
rect 128556 336776 129646 336832
rect 129702 336776 129707 336832
rect 128556 336774 129707 336776
rect 128556 336772 128562 336774
rect 129641 336771 129707 336774
rect 364517 336834 364583 336837
rect 371233 336836 371299 336837
rect 365478 336834 365484 336836
rect 364517 336832 365484 336834
rect 364517 336776 364522 336832
rect 364578 336776 365484 336832
rect 364517 336774 365484 336776
rect 364517 336771 364583 336774
rect 365478 336772 365484 336774
rect 365548 336772 365554 336836
rect 371182 336772 371188 336836
rect 371252 336834 371299 336836
rect 376845 336836 376911 336837
rect 376845 336834 376892 336836
rect 371252 336832 371344 336834
rect 371294 336776 371344 336832
rect 371252 336774 371344 336776
rect 376800 336832 376892 336834
rect 376800 336776 376850 336832
rect 376800 336774 376892 336776
rect 371252 336772 371299 336774
rect 371233 336771 371299 336772
rect 376845 336772 376892 336774
rect 376956 336772 376962 336836
rect 390553 336834 390619 336837
rect 391238 336834 391244 336836
rect 390553 336832 391244 336834
rect 390553 336776 390558 336832
rect 390614 336776 391244 336832
rect 390553 336774 391244 336776
rect 376845 336771 376911 336772
rect 390553 336771 390619 336774
rect 391238 336772 391244 336774
rect 391308 336772 391314 336836
rect 397453 336834 397519 336837
rect 398414 336834 398420 336836
rect 397453 336832 398420 336834
rect 397453 336776 397458 336832
rect 397514 336776 398420 336832
rect 397453 336774 398420 336776
rect 397453 336771 397519 336774
rect 398414 336772 398420 336774
rect 398484 336772 398490 336836
rect 403249 336834 403315 336837
rect 403566 336834 403572 336836
rect 403249 336832 403572 336834
rect 403249 336776 403254 336832
rect 403310 336776 403572 336832
rect 403249 336774 403572 336776
rect 403249 336771 403315 336774
rect 403566 336772 403572 336774
rect 403636 336772 403642 336836
rect -960 332196 480 332436
rect 579981 325274 580047 325277
rect 583520 325274 584960 325364
rect 579981 325272 584960 325274
rect 579981 325216 579986 325272
rect 580042 325216 584960 325272
rect 579981 325214 584960 325216
rect 579981 325211 580047 325214
rect 583520 325124 584960 325214
rect -960 319290 480 319380
rect 3417 319290 3483 319293
rect -960 319288 3483 319290
rect -960 319232 3422 319288
rect 3478 319232 3483 319288
rect -960 319230 3483 319232
rect -960 319140 480 319230
rect 3417 319227 3483 319230
rect 580165 312082 580231 312085
rect 583520 312082 584960 312172
rect 580165 312080 584960 312082
rect 580165 312024 580170 312080
rect 580226 312024 584960 312080
rect 580165 312022 584960 312024
rect 580165 312019 580231 312022
rect 583520 311932 584960 312022
rect -960 306234 480 306324
rect 3417 306234 3483 306237
rect -960 306232 3483 306234
rect -960 306176 3422 306232
rect 3478 306176 3483 306232
rect -960 306174 3483 306176
rect -960 306084 480 306174
rect 3417 306171 3483 306174
rect 580165 298754 580231 298757
rect 583520 298754 584960 298844
rect 580165 298752 584960 298754
rect 580165 298696 580170 298752
rect 580226 298696 584960 298752
rect 580165 298694 584960 298696
rect 580165 298691 580231 298694
rect 583520 298604 584960 298694
rect -960 293178 480 293268
rect 3417 293178 3483 293181
rect -960 293176 3483 293178
rect -960 293120 3422 293176
rect 3478 293120 3483 293176
rect -960 293118 3483 293120
rect -960 293028 480 293118
rect 3417 293115 3483 293118
rect 583520 285276 584960 285516
rect -960 279972 480 280212
rect 580165 272234 580231 272237
rect 583520 272234 584960 272324
rect 580165 272232 584960 272234
rect 580165 272176 580170 272232
rect 580226 272176 584960 272232
rect 580165 272174 584960 272176
rect 580165 272171 580231 272174
rect 583520 272084 584960 272174
rect -960 267202 480 267292
rect 3049 267202 3115 267205
rect -960 267200 3115 267202
rect -960 267144 3054 267200
rect 3110 267144 3115 267200
rect -960 267142 3115 267144
rect -960 267052 480 267142
rect 3049 267139 3115 267142
rect 580165 258906 580231 258909
rect 583520 258906 584960 258996
rect 580165 258904 584960 258906
rect 580165 258848 580170 258904
rect 580226 258848 584960 258904
rect 580165 258846 584960 258848
rect 580165 258843 580231 258846
rect 583520 258756 584960 258846
rect -960 254146 480 254236
rect 3417 254146 3483 254149
rect -960 254144 3483 254146
rect -960 254088 3422 254144
rect 3478 254088 3483 254144
rect -960 254086 3483 254088
rect -960 253996 480 254086
rect 3417 254083 3483 254086
rect 579613 245578 579679 245581
rect 583520 245578 584960 245668
rect 579613 245576 584960 245578
rect 579613 245520 579618 245576
rect 579674 245520 584960 245576
rect 579613 245518 584960 245520
rect 579613 245515 579679 245518
rect 583520 245428 584960 245518
rect 40585 242994 40651 242997
rect 265617 242994 265683 242997
rect 40585 242992 265683 242994
rect 40585 242936 40590 242992
rect 40646 242936 265622 242992
rect 265678 242936 265683 242992
rect 40585 242934 265683 242936
rect 40585 242931 40651 242934
rect 265617 242931 265683 242934
rect 43069 241634 43135 241637
rect 168465 241634 168531 241637
rect 43069 241632 168531 241634
rect 43069 241576 43074 241632
rect 43130 241576 168470 241632
rect 168526 241576 168531 241632
rect 43069 241574 168531 241576
rect 43069 241571 43135 241574
rect 168465 241571 168531 241574
rect -960 241090 480 241180
rect 3417 241090 3483 241093
rect -960 241088 3483 241090
rect -960 241032 3422 241088
rect 3478 241032 3483 241088
rect -960 241030 3483 241032
rect -960 240940 480 241030
rect 3417 241027 3483 241030
rect 45921 239866 45987 239869
rect 73429 239868 73495 239869
rect 73429 239866 73476 239868
rect 45921 239864 55230 239866
rect 45921 239808 45926 239864
rect 45982 239808 55230 239864
rect 45921 239806 55230 239808
rect 73384 239864 73476 239866
rect 73384 239808 73434 239864
rect 73384 239806 73476 239808
rect 45921 239803 45987 239806
rect 50981 239730 51047 239733
rect 50981 239728 53114 239730
rect 50981 239672 50986 239728
rect 51042 239672 53114 239728
rect 50981 239670 53114 239672
rect 50981 239667 51047 239670
rect 53054 238778 53114 239670
rect 55170 238914 55230 239806
rect 73429 239804 73476 239806
rect 73540 239804 73546 239868
rect 73429 239803 73495 239804
rect 57697 239732 57763 239733
rect 59169 239732 59235 239733
rect 57646 239730 57652 239732
rect 57606 239670 57652 239730
rect 57716 239728 57763 239732
rect 59118 239730 59124 239732
rect 57758 239672 57763 239728
rect 57646 239668 57652 239670
rect 57716 239668 57763 239672
rect 59078 239670 59124 239730
rect 59188 239728 59235 239732
rect 75821 239732 75887 239733
rect 75821 239730 75868 239732
rect 59230 239672 59235 239728
rect 59118 239668 59124 239670
rect 59188 239668 59235 239672
rect 75776 239728 75868 239730
rect 75776 239672 75826 239728
rect 75776 239670 75868 239672
rect 57697 239667 57763 239668
rect 59169 239667 59235 239668
rect 75821 239668 75868 239670
rect 75932 239668 75938 239732
rect 87137 239730 87203 239733
rect 84150 239728 87203 239730
rect 84150 239672 87142 239728
rect 87198 239672 87203 239728
rect 84150 239670 87203 239672
rect 75821 239667 75887 239668
rect 59302 239396 59308 239460
rect 59372 239458 59378 239460
rect 84150 239458 84210 239670
rect 87137 239667 87203 239670
rect 59372 239398 84210 239458
rect 59372 239396 59378 239398
rect 276657 238914 276723 238917
rect 55170 238912 276723 238914
rect 55170 238856 276662 238912
rect 276718 238856 276723 238912
rect 55170 238854 276723 238856
rect 276657 238851 276723 238854
rect 283557 238778 283623 238781
rect 53054 238776 283623 238778
rect 53054 238720 283562 238776
rect 283618 238720 283623 238776
rect 53054 238718 283623 238720
rect 283557 238715 283623 238718
rect 40125 238098 40191 238101
rect 40125 238096 40234 238098
rect 40125 238040 40130 238096
rect 40186 238040 40234 238096
rect 40125 238035 40234 238040
rect 40174 237524 40234 238035
rect 241145 237826 241211 237829
rect 238004 237824 241211 237826
rect 238004 237768 241150 237824
rect 241206 237768 241211 237824
rect 238004 237766 241211 237768
rect 241145 237763 241211 237766
rect 240593 232794 240659 232797
rect 238004 232792 240659 232794
rect 238004 232736 240598 232792
rect 240654 232736 240659 232792
rect 238004 232734 240659 232736
rect 240593 232731 240659 232734
rect 580717 232386 580783 232389
rect 583520 232386 584960 232476
rect 580717 232384 584960 232386
rect 580717 232328 580722 232384
rect 580778 232328 584960 232384
rect 580717 232326 584960 232328
rect 580717 232323 580783 232326
rect 583520 232236 584960 232326
rect 38561 232114 38627 232117
rect 38561 232112 40204 232114
rect 38561 232056 38566 232112
rect 38622 232056 40204 232112
rect 38561 232054 40204 232056
rect 38561 232051 38627 232054
rect -960 227884 480 228124
rect 240133 227762 240199 227765
rect 238004 227760 240199 227762
rect 238004 227704 240138 227760
rect 240194 227704 240199 227760
rect 238004 227702 240199 227704
rect 240133 227699 240199 227702
rect 39481 226674 39547 226677
rect 39481 226672 40204 226674
rect 39481 226616 39486 226672
rect 39542 226616 40204 226672
rect 39481 226614 40204 226616
rect 39481 226611 39547 226614
rect 240869 222730 240935 222733
rect 238004 222728 240935 222730
rect 238004 222672 240874 222728
rect 240930 222672 240935 222728
rect 238004 222670 240935 222672
rect 240869 222667 240935 222670
rect 39389 221234 39455 221237
rect 39389 221232 40204 221234
rect 39389 221176 39394 221232
rect 39450 221176 40204 221232
rect 39389 221174 40204 221176
rect 39389 221171 39455 221174
rect 580625 219058 580691 219061
rect 583520 219058 584960 219148
rect 580625 219056 584960 219058
rect 580625 219000 580630 219056
rect 580686 219000 584960 219056
rect 580625 218998 584960 219000
rect 580625 218995 580691 218998
rect 583520 218908 584960 218998
rect 239489 217698 239555 217701
rect 238004 217696 239555 217698
rect 238004 217640 239494 217696
rect 239550 217640 239555 217696
rect 238004 217638 239555 217640
rect 239489 217635 239555 217638
rect 36537 215794 36603 215797
rect 36537 215792 40204 215794
rect 36537 215736 36542 215792
rect 36598 215736 40204 215792
rect 36537 215734 40204 215736
rect 36537 215731 36603 215734
rect -960 214978 480 215068
rect 3325 214978 3391 214981
rect -960 214976 3391 214978
rect -960 214920 3330 214976
rect 3386 214920 3391 214976
rect -960 214918 3391 214920
rect -960 214828 480 214918
rect 3325 214915 3391 214918
rect 241237 212802 241303 212805
rect 238004 212800 241303 212802
rect 238004 212744 241242 212800
rect 241298 212744 241303 212800
rect 238004 212742 241303 212744
rect 241237 212739 241303 212742
rect 36629 210490 36695 210493
rect 36629 210488 40204 210490
rect 36629 210432 36634 210488
rect 36690 210432 40204 210488
rect 36629 210430 40204 210432
rect 36629 210427 36695 210430
rect 241421 207770 241487 207773
rect 238004 207768 241487 207770
rect 238004 207712 241426 207768
rect 241482 207712 241487 207768
rect 238004 207710 241487 207712
rect 241421 207707 241487 207710
rect 579797 205730 579863 205733
rect 583520 205730 584960 205820
rect 579797 205728 584960 205730
rect 579797 205672 579802 205728
rect 579858 205672 584960 205728
rect 579797 205670 584960 205672
rect 579797 205667 579863 205670
rect 583520 205580 584960 205670
rect 39205 205050 39271 205053
rect 39205 205048 40204 205050
rect 39205 204992 39210 205048
rect 39266 204992 40204 205048
rect 39205 204990 40204 204992
rect 39205 204987 39271 204990
rect 241421 202738 241487 202741
rect 238004 202736 241487 202738
rect 238004 202680 241426 202736
rect 241482 202680 241487 202736
rect 238004 202678 241487 202680
rect 241421 202675 241487 202678
rect -960 201922 480 202012
rect 3049 201922 3115 201925
rect -960 201920 3115 201922
rect -960 201864 3054 201920
rect 3110 201864 3115 201920
rect -960 201862 3115 201864
rect -960 201772 480 201862
rect 3049 201859 3115 201862
rect 37733 199610 37799 199613
rect 37733 199608 40204 199610
rect 37733 199552 37738 199608
rect 37794 199552 40204 199608
rect 37733 199550 40204 199552
rect 37733 199547 37799 199550
rect 241421 197706 241487 197709
rect 238004 197704 241487 197706
rect 238004 197648 241426 197704
rect 241482 197648 241487 197704
rect 238004 197646 241487 197648
rect 241421 197643 241487 197646
rect 39113 194170 39179 194173
rect 39113 194168 40204 194170
rect 39113 194112 39118 194168
rect 39174 194112 40204 194168
rect 39113 194110 40204 194112
rect 39113 194107 39179 194110
rect 240593 192674 240659 192677
rect 238004 192672 240659 192674
rect 238004 192616 240598 192672
rect 240654 192616 240659 192672
rect 238004 192614 240659 192616
rect 240593 192611 240659 192614
rect 579613 192538 579679 192541
rect 583520 192538 584960 192628
rect 579613 192536 584960 192538
rect 579613 192480 579618 192536
rect 579674 192480 584960 192536
rect 579613 192478 584960 192480
rect 579613 192475 579679 192478
rect 583520 192388 584960 192478
rect -960 188866 480 188956
rect 3509 188866 3575 188869
rect -960 188864 3575 188866
rect -960 188808 3514 188864
rect 3570 188808 3575 188864
rect -960 188806 3575 188808
rect -960 188716 480 188806
rect 3509 188803 3575 188806
rect 37825 188730 37891 188733
rect 37825 188728 40204 188730
rect 37825 188672 37830 188728
rect 37886 188672 40204 188728
rect 37825 188670 40204 188672
rect 37825 188667 37891 188670
rect 241421 187642 241487 187645
rect 238004 187640 241487 187642
rect 238004 187584 241426 187640
rect 241482 187584 241487 187640
rect 238004 187582 241487 187584
rect 241421 187579 241487 187582
rect 36813 183426 36879 183429
rect 36813 183424 40204 183426
rect 36813 183368 36818 183424
rect 36874 183368 40204 183424
rect 36813 183366 40204 183368
rect 36813 183363 36879 183366
rect 241421 182746 241487 182749
rect 238004 182744 241487 182746
rect 238004 182688 241426 182744
rect 241482 182688 241487 182744
rect 238004 182686 241487 182688
rect 241421 182683 241487 182686
rect 580533 179210 580599 179213
rect 583520 179210 584960 179300
rect 580533 179208 584960 179210
rect 580533 179152 580538 179208
rect 580594 179152 584960 179208
rect 580533 179150 584960 179152
rect 580533 179147 580599 179150
rect 583520 179060 584960 179150
rect 36721 177986 36787 177989
rect 36721 177984 40204 177986
rect 36721 177928 36726 177984
rect 36782 177928 40204 177984
rect 36721 177926 40204 177928
rect 36721 177923 36787 177926
rect 240133 177714 240199 177717
rect 238004 177712 240199 177714
rect 238004 177656 240138 177712
rect 240194 177656 240199 177712
rect 238004 177654 240199 177656
rect 240133 177651 240199 177654
rect -960 175796 480 176036
rect 241237 172682 241303 172685
rect 238004 172680 241303 172682
rect 238004 172624 241242 172680
rect 241298 172624 241303 172680
rect 238004 172622 241303 172624
rect 241237 172619 241303 172622
rect 38745 172546 38811 172549
rect 38745 172544 40204 172546
rect 38745 172488 38750 172544
rect 38806 172488 40204 172544
rect 38745 172486 40204 172488
rect 38745 172483 38811 172486
rect 239305 167650 239371 167653
rect 238004 167648 239371 167650
rect 238004 167592 239310 167648
rect 239366 167592 239371 167648
rect 238004 167590 239371 167592
rect 239305 167587 239371 167590
rect 37917 167106 37983 167109
rect 37917 167104 40204 167106
rect 37917 167048 37922 167104
rect 37978 167048 40204 167104
rect 37917 167046 40204 167048
rect 37917 167043 37983 167046
rect 580165 165882 580231 165885
rect 583520 165882 584960 165972
rect 580165 165880 584960 165882
rect 580165 165824 580170 165880
rect 580226 165824 584960 165880
rect 580165 165822 584960 165824
rect 580165 165819 580231 165822
rect 583520 165732 584960 165822
rect -960 162890 480 162980
rect 3233 162890 3299 162893
rect -960 162888 3299 162890
rect -960 162832 3238 162888
rect 3294 162832 3299 162888
rect -960 162830 3299 162832
rect -960 162740 480 162830
rect 3233 162827 3299 162830
rect 237974 162346 238034 162588
rect 238109 162346 238175 162349
rect 237974 162344 238175 162346
rect 237974 162288 238114 162344
rect 238170 162288 238175 162344
rect 237974 162286 238175 162288
rect 238109 162283 238175 162286
rect 36905 161666 36971 161669
rect 36905 161664 40204 161666
rect 36905 161608 36910 161664
rect 36966 161608 40204 161664
rect 36905 161606 40204 161608
rect 36905 161603 36971 161606
rect 241053 157586 241119 157589
rect 238004 157584 241119 157586
rect 238004 157528 241058 157584
rect 241114 157528 241119 157584
rect 238004 157526 241119 157528
rect 241053 157523 241119 157526
rect 38009 156362 38075 156365
rect 38009 156360 40204 156362
rect 38009 156304 38014 156360
rect 38070 156304 40204 156360
rect 38009 156302 40204 156304
rect 38009 156299 38075 156302
rect 240501 152690 240567 152693
rect 238004 152688 240567 152690
rect 238004 152632 240506 152688
rect 240562 152632 240567 152688
rect 238004 152630 240567 152632
rect 240501 152627 240567 152630
rect 580441 152690 580507 152693
rect 583520 152690 584960 152780
rect 580441 152688 584960 152690
rect 580441 152632 580446 152688
rect 580502 152632 584960 152688
rect 580441 152630 584960 152632
rect 580441 152627 580507 152630
rect 583520 152540 584960 152630
rect 37733 150922 37799 150925
rect 37733 150920 40204 150922
rect 37733 150864 37738 150920
rect 37794 150864 40204 150920
rect 37733 150862 40204 150864
rect 37733 150859 37799 150862
rect -960 149834 480 149924
rect 3509 149834 3575 149837
rect -960 149832 3575 149834
rect -960 149776 3514 149832
rect 3570 149776 3575 149832
rect -960 149774 3575 149776
rect -960 149684 480 149774
rect 3509 149771 3575 149774
rect 239213 147658 239279 147661
rect 238004 147656 239279 147658
rect 238004 147600 239218 147656
rect 239274 147600 239279 147656
rect 238004 147598 239279 147600
rect 239213 147595 239279 147598
rect 37089 145482 37155 145485
rect 37089 145480 40204 145482
rect 37089 145424 37094 145480
rect 37150 145424 40204 145480
rect 37089 145422 40204 145424
rect 37089 145419 37155 145422
rect 241145 142626 241211 142629
rect 238004 142624 241211 142626
rect 238004 142568 241150 142624
rect 241206 142568 241211 142624
rect 238004 142566 241211 142568
rect 241145 142563 241211 142566
rect 39021 140042 39087 140045
rect 39021 140040 40204 140042
rect 39021 139984 39026 140040
rect 39082 139984 40204 140040
rect 39021 139982 40204 139984
rect 39021 139979 39087 139982
rect 580165 139362 580231 139365
rect 583520 139362 584960 139452
rect 580165 139360 584960 139362
rect 580165 139304 580170 139360
rect 580226 139304 584960 139360
rect 580165 139302 584960 139304
rect 580165 139299 580231 139302
rect 583520 139212 584960 139302
rect 241421 137594 241487 137597
rect 238004 137592 241487 137594
rect 238004 137536 241426 137592
rect 241482 137536 241487 137592
rect 238004 137534 241487 137536
rect 241421 137531 241487 137534
rect -960 136778 480 136868
rect 3509 136778 3575 136781
rect -960 136776 3575 136778
rect -960 136720 3514 136776
rect 3570 136720 3575 136776
rect -960 136718 3575 136720
rect -960 136628 480 136718
rect 3509 136715 3575 136718
rect 38009 134602 38075 134605
rect 38009 134600 40204 134602
rect 38009 134544 38014 134600
rect 38070 134544 40204 134600
rect 38009 134542 40204 134544
rect 38009 134539 38075 134542
rect 240685 132562 240751 132565
rect 238004 132560 240751 132562
rect 238004 132504 240690 132560
rect 240746 132504 240751 132560
rect 238004 132502 240751 132504
rect 240685 132499 240751 132502
rect 37549 129162 37615 129165
rect 37549 129160 40204 129162
rect 37549 129104 37554 129160
rect 37610 129104 40204 129160
rect 37549 129102 40204 129104
rect 37549 129099 37615 129102
rect 241421 127666 241487 127669
rect 238004 127664 241487 127666
rect 238004 127608 241426 127664
rect 241482 127608 241487 127664
rect 238004 127606 241487 127608
rect 241421 127603 241487 127606
rect 580165 126034 580231 126037
rect 583520 126034 584960 126124
rect 580165 126032 584960 126034
rect 580165 125976 580170 126032
rect 580226 125976 584960 126032
rect 580165 125974 584960 125976
rect 580165 125971 580231 125974
rect 583520 125884 584960 125974
rect 38009 123858 38075 123861
rect 38009 123856 40204 123858
rect -960 123572 480 123812
rect 38009 123800 38014 123856
rect 38070 123800 40204 123856
rect 38009 123798 40204 123800
rect 38009 123795 38075 123798
rect 238753 122634 238819 122637
rect 238004 122632 238819 122634
rect 238004 122576 238758 122632
rect 238814 122576 238819 122632
rect 238004 122574 238819 122576
rect 238753 122571 238819 122574
rect 38929 118418 38995 118421
rect 38929 118416 40204 118418
rect 38929 118360 38934 118416
rect 38990 118360 40204 118416
rect 38929 118358 40204 118360
rect 38929 118355 38995 118358
rect 241697 117602 241763 117605
rect 238004 117600 241763 117602
rect 238004 117544 241702 117600
rect 241758 117544 241763 117600
rect 238004 117542 241763 117544
rect 241697 117539 241763 117542
rect 38101 112978 38167 112981
rect 38101 112976 40204 112978
rect 38101 112920 38106 112976
rect 38162 112920 40204 112976
rect 38101 112918 40204 112920
rect 38101 112915 38167 112918
rect 579613 112842 579679 112845
rect 583520 112842 584960 112932
rect 579613 112840 584960 112842
rect 579613 112784 579618 112840
rect 579674 112784 584960 112840
rect 579613 112782 584960 112784
rect 579613 112779 579679 112782
rect 583520 112692 584960 112782
rect 240869 112570 240935 112573
rect 238004 112568 240935 112570
rect 238004 112512 240874 112568
rect 240930 112512 240935 112568
rect 238004 112510 240935 112512
rect 240869 112507 240935 112510
rect -960 110666 480 110756
rect 3141 110666 3207 110669
rect -960 110664 3207 110666
rect -960 110608 3146 110664
rect 3202 110608 3207 110664
rect -960 110606 3207 110608
rect -960 110516 480 110606
rect 3141 110603 3207 110606
rect 38009 107538 38075 107541
rect 241421 107538 241487 107541
rect 38009 107536 40204 107538
rect 38009 107480 38014 107536
rect 38070 107480 40204 107536
rect 38009 107478 40204 107480
rect 238004 107536 241487 107538
rect 238004 107480 241426 107536
rect 241482 107480 241487 107536
rect 238004 107478 241487 107480
rect 38009 107475 38075 107478
rect 241421 107475 241487 107478
rect 241237 102506 241303 102509
rect 238004 102504 241303 102506
rect 238004 102448 241242 102504
rect 241298 102448 241303 102504
rect 238004 102446 241303 102448
rect 241237 102443 241303 102446
rect 37825 102098 37891 102101
rect 37825 102096 40204 102098
rect 37825 102040 37830 102096
rect 37886 102040 40204 102096
rect 37825 102038 40204 102040
rect 37825 102035 37891 102038
rect 580165 99514 580231 99517
rect 583520 99514 584960 99604
rect 580165 99512 584960 99514
rect 580165 99456 580170 99512
rect 580226 99456 584960 99512
rect 580165 99454 584960 99456
rect 580165 99451 580231 99454
rect 583520 99364 584960 99454
rect -960 97610 480 97700
rect 3417 97610 3483 97613
rect 239121 97610 239187 97613
rect -960 97608 3483 97610
rect -960 97552 3422 97608
rect 3478 97552 3483 97608
rect -960 97550 3483 97552
rect 238004 97608 239187 97610
rect 238004 97552 239126 97608
rect 239182 97552 239187 97608
rect 238004 97550 239187 97552
rect -960 97460 480 97550
rect 3417 97547 3483 97550
rect 239121 97547 239187 97550
rect 38285 96794 38351 96797
rect 38285 96792 40204 96794
rect 38285 96736 38290 96792
rect 38346 96736 40204 96792
rect 38285 96734 40204 96736
rect 38285 96731 38351 96734
rect 241421 92578 241487 92581
rect 238004 92576 241487 92578
rect 238004 92520 241426 92576
rect 241482 92520 241487 92576
rect 238004 92518 241487 92520
rect 241421 92515 241487 92518
rect 38837 91354 38903 91357
rect 38837 91352 40204 91354
rect 38837 91296 38842 91352
rect 38898 91296 40204 91352
rect 38837 91294 40204 91296
rect 38837 91291 38903 91294
rect 241421 87546 241487 87549
rect 238004 87544 241487 87546
rect 238004 87488 241426 87544
rect 241482 87488 241487 87544
rect 238004 87486 241487 87488
rect 241421 87483 241487 87486
rect 579613 86186 579679 86189
rect 583520 86186 584960 86276
rect 579613 86184 584960 86186
rect 579613 86128 579618 86184
rect 579674 86128 584960 86184
rect 579613 86126 584960 86128
rect 579613 86123 579679 86126
rect 583520 86036 584960 86126
rect 37181 85914 37247 85917
rect 37181 85912 40204 85914
rect 37181 85856 37186 85912
rect 37242 85856 40204 85912
rect 37181 85854 40204 85856
rect 37181 85851 37247 85854
rect -960 84690 480 84780
rect 3141 84690 3207 84693
rect -960 84688 3207 84690
rect -960 84632 3146 84688
rect 3202 84632 3207 84688
rect -960 84630 3207 84632
rect -960 84540 480 84630
rect 3141 84627 3207 84630
rect 240317 82514 240383 82517
rect 238004 82512 240383 82514
rect 238004 82456 240322 82512
rect 240378 82456 240383 82512
rect 238004 82454 240383 82456
rect 240317 82451 240383 82454
rect 38377 80474 38443 80477
rect 38377 80472 40204 80474
rect 38377 80416 38382 80472
rect 38438 80416 40204 80472
rect 38377 80414 40204 80416
rect 38377 80411 38443 80414
rect 241237 77482 241303 77485
rect 238004 77480 241303 77482
rect 238004 77424 241242 77480
rect 241298 77424 241303 77480
rect 238004 77422 241303 77424
rect 241237 77419 241303 77422
rect 38009 75034 38075 75037
rect 38009 75032 40204 75034
rect 38009 74976 38014 75032
rect 38070 74976 40204 75032
rect 38009 74974 40204 74976
rect 38009 74971 38075 74974
rect 580165 72994 580231 72997
rect 583520 72994 584960 73084
rect 580165 72992 584960 72994
rect 580165 72936 580170 72992
rect 580226 72936 584960 72992
rect 580165 72934 584960 72936
rect 580165 72931 580231 72934
rect 583520 72844 584960 72934
rect 240409 72450 240475 72453
rect 238004 72448 240475 72450
rect 238004 72392 240414 72448
rect 240470 72392 240475 72448
rect 238004 72390 240475 72392
rect 240409 72387 240475 72390
rect -960 71634 480 71724
rect 3141 71634 3207 71637
rect -960 71632 3207 71634
rect -960 71576 3146 71632
rect 3202 71576 3207 71632
rect -960 71574 3207 71576
rect -960 71484 480 71574
rect 3141 71571 3207 71574
rect 38561 69730 38627 69733
rect 38561 69728 40204 69730
rect 38561 69672 38566 69728
rect 38622 69672 40204 69728
rect 38561 69670 40204 69672
rect 38561 69667 38627 69670
rect 241421 67554 241487 67557
rect 238004 67552 241487 67554
rect 238004 67496 241426 67552
rect 241482 67496 241487 67552
rect 238004 67494 241487 67496
rect 241421 67491 241487 67494
rect 38193 64290 38259 64293
rect 38193 64288 40204 64290
rect 38193 64232 38198 64288
rect 38254 64232 40204 64288
rect 38193 64230 40204 64232
rect 38193 64227 38259 64230
rect 241237 62522 241303 62525
rect 238004 62520 241303 62522
rect 238004 62464 241242 62520
rect 241298 62464 241303 62520
rect 238004 62462 241303 62464
rect 241237 62459 241303 62462
rect 580349 59666 580415 59669
rect 583520 59666 584960 59756
rect 580349 59664 584960 59666
rect 580349 59608 580354 59664
rect 580410 59608 584960 59664
rect 580349 59606 584960 59608
rect 580349 59603 580415 59606
rect 583520 59516 584960 59606
rect 38653 58850 38719 58853
rect 38653 58848 40204 58850
rect 38653 58792 38658 58848
rect 38714 58792 40204 58848
rect 38653 58790 40204 58792
rect 38653 58787 38719 58790
rect -960 58578 480 58668
rect 3049 58578 3115 58581
rect -960 58576 3115 58578
rect -960 58520 3054 58576
rect 3110 58520 3115 58576
rect -960 58518 3115 58520
rect -960 58428 480 58518
rect 3049 58515 3115 58518
rect 237925 57898 237991 57901
rect 237925 57896 238034 57898
rect 237925 57840 237930 57896
rect 237986 57840 238034 57896
rect 237925 57835 238034 57840
rect 237974 57460 238034 57835
rect 36997 53410 37063 53413
rect 36997 53408 40204 53410
rect 36997 53352 37002 53408
rect 37058 53352 40204 53408
rect 36997 53350 40204 53352
rect 36997 53347 37063 53350
rect 241421 52458 241487 52461
rect 238004 52456 241487 52458
rect 238004 52400 241426 52456
rect 241482 52400 241487 52456
rect 238004 52398 241487 52400
rect 241421 52395 241487 52398
rect 40542 47428 40602 47940
rect 40534 47364 40540 47428
rect 40604 47364 40610 47428
rect 240225 47426 240291 47429
rect 238004 47424 240291 47426
rect 238004 47368 240230 47424
rect 240286 47368 240291 47424
rect 238004 47366 240291 47368
rect 240225 47363 240291 47366
rect 580165 46338 580231 46341
rect 583520 46338 584960 46428
rect 580165 46336 584960 46338
rect 580165 46280 580170 46336
rect 580226 46280 584960 46336
rect 580165 46278 584960 46280
rect 580165 46275 580231 46278
rect 583520 46188 584960 46278
rect -960 45522 480 45612
rect 3417 45522 3483 45525
rect -960 45520 3483 45522
rect -960 45464 3422 45520
rect 3478 45464 3483 45520
rect -960 45462 3483 45464
rect -960 45372 480 45462
rect 3417 45459 3483 45462
rect 38561 45522 38627 45525
rect 40534 45522 40540 45524
rect 38561 45520 40540 45522
rect 38561 45464 38566 45520
rect 38622 45464 40540 45520
rect 38561 45462 40540 45464
rect 38561 45459 38627 45462
rect 40534 45460 40540 45462
rect 40604 45460 40610 45524
rect 38009 42666 38075 42669
rect 38009 42664 40204 42666
rect 38009 42608 38014 42664
rect 38070 42608 40204 42664
rect 38009 42606 40204 42608
rect 38009 42603 38075 42606
rect 238937 42530 239003 42533
rect 238004 42528 239003 42530
rect 238004 42472 238942 42528
rect 238998 42472 239003 42528
rect 238004 42470 239003 42472
rect 238937 42467 239003 42470
rect 237557 41170 237623 41173
rect 238201 41170 238267 41173
rect 237557 41168 238267 41170
rect 237557 41112 237562 41168
rect 237618 41112 238206 41168
rect 238262 41112 238267 41168
rect 237557 41110 238267 41112
rect 237557 41107 237623 41110
rect 238201 41107 238267 41110
rect 237741 41034 237807 41037
rect 238109 41034 238175 41037
rect 237741 41032 238175 41034
rect 237741 40976 237746 41032
rect 237802 40976 238114 41032
rect 238170 40976 238175 41032
rect 237741 40974 238175 40976
rect 237741 40971 237807 40974
rect 238109 40971 238175 40974
rect 237649 40898 237715 40901
rect 237925 40898 237991 40901
rect 237649 40896 237991 40898
rect 237649 40840 237654 40896
rect 237710 40840 237930 40896
rect 237986 40840 237991 40896
rect 237649 40838 237991 40840
rect 237649 40835 237715 40838
rect 237925 40835 237991 40838
rect 58249 39948 58315 39949
rect 58198 39946 58204 39948
rect 58158 39886 58204 39946
rect 58268 39944 58315 39948
rect 58310 39888 58315 39944
rect 58198 39884 58204 39886
rect 58268 39884 58315 39888
rect 58249 39883 58315 39884
rect 52310 38524 52316 38588
rect 52380 38586 52386 38588
rect 203333 38586 203399 38589
rect 52380 38584 203399 38586
rect 52380 38528 203338 38584
rect 203394 38528 203399 38584
rect 52380 38526 203399 38528
rect 52380 38524 52386 38526
rect 203333 38523 203399 38526
rect 215201 38586 215267 38589
rect 233182 38586 233188 38588
rect 215201 38584 233188 38586
rect 215201 38528 215206 38584
rect 215262 38528 233188 38584
rect 215201 38526 233188 38528
rect 215201 38523 215267 38526
rect 233182 38524 233188 38526
rect 233252 38524 233258 38588
rect 57646 38388 57652 38452
rect 57716 38450 57722 38452
rect 207289 38450 207355 38453
rect 57716 38448 207355 38450
rect 57716 38392 207294 38448
rect 207350 38392 207355 38448
rect 57716 38390 207355 38392
rect 57716 38388 57722 38390
rect 207289 38387 207355 38390
rect 216489 38450 216555 38453
rect 231894 38450 231900 38452
rect 216489 38448 231900 38450
rect 216489 38392 216494 38448
rect 216550 38392 231900 38448
rect 216489 38390 231900 38392
rect 216489 38387 216555 38390
rect 231894 38388 231900 38390
rect 231964 38388 231970 38452
rect 59118 38252 59124 38316
rect 59188 38314 59194 38316
rect 204713 38314 204779 38317
rect 59188 38312 204779 38314
rect 59188 38256 204718 38312
rect 204774 38256 204779 38312
rect 59188 38254 204779 38256
rect 59188 38252 59194 38254
rect 204713 38251 204779 38254
rect 59302 38116 59308 38180
rect 59372 38178 59378 38180
rect 200757 38178 200823 38181
rect 59372 38176 200823 38178
rect 59372 38120 200762 38176
rect 200818 38120 200823 38176
rect 59372 38118 200823 38120
rect 59372 38116 59378 38118
rect 200757 38115 200823 38118
rect 56358 37980 56364 38044
rect 56428 38042 56434 38044
rect 192845 38042 192911 38045
rect 56428 38040 192911 38042
rect 56428 37984 192850 38040
rect 192906 37984 192911 38040
rect 56428 37982 192911 37984
rect 56428 37980 56434 37982
rect 192845 37979 192911 37982
rect 53598 37844 53604 37908
rect 53668 37906 53674 37908
rect 188889 37906 188955 37909
rect 53668 37904 188955 37906
rect 53668 37848 188894 37904
rect 188950 37848 188955 37904
rect 53668 37846 188955 37848
rect 53668 37844 53674 37846
rect 188889 37843 188955 37846
rect 57830 37708 57836 37772
rect 57900 37770 57906 37772
rect 187601 37770 187667 37773
rect 57900 37768 187667 37770
rect 57900 37712 187606 37768
rect 187662 37712 187667 37768
rect 57900 37710 187667 37712
rect 57900 37708 57906 37710
rect 187601 37707 187667 37710
rect 580165 33146 580231 33149
rect 583520 33146 584960 33236
rect 580165 33144 584960 33146
rect 580165 33088 580170 33144
rect 580226 33088 584960 33144
rect 580165 33086 584960 33088
rect 580165 33083 580231 33086
rect 583520 32996 584960 33086
rect -960 32466 480 32556
rect 2865 32466 2931 32469
rect -960 32464 2931 32466
rect -960 32408 2870 32464
rect 2926 32408 2931 32464
rect -960 32406 2931 32408
rect -960 32316 480 32406
rect 2865 32403 2931 32406
rect 580257 19818 580323 19821
rect 583520 19818 584960 19908
rect 580257 19816 584960 19818
rect 580257 19760 580262 19816
rect 580318 19760 584960 19816
rect 580257 19758 584960 19760
rect 580257 19755 580323 19758
rect 583520 19668 584960 19758
rect -960 19410 480 19500
rect 3417 19410 3483 19413
rect -960 19408 3483 19410
rect -960 19352 3422 19408
rect 3478 19352 3483 19408
rect -960 19350 3483 19352
rect -960 19260 480 19350
rect 3417 19347 3483 19350
rect 580165 6626 580231 6629
rect 583520 6626 584960 6716
rect 580165 6624 584960 6626
rect -960 6490 480 6580
rect 580165 6568 580170 6624
rect 580226 6568 584960 6624
rect 580165 6566 584960 6568
rect 580165 6563 580231 6566
rect 3417 6490 3483 6493
rect -960 6488 3483 6490
rect -960 6432 3422 6488
rect 3478 6432 3483 6488
rect 583520 6476 584960 6566
rect -960 6430 3483 6432
rect -960 6340 480 6430
rect 3417 6427 3483 6430
<< via3 >>
rect 76972 338132 77036 338196
rect 80652 338132 80716 338196
rect 83964 338132 84028 338196
rect 90956 338132 91020 338196
rect 98500 338132 98564 338196
rect 131068 338132 131132 338196
rect 372292 338132 372356 338196
rect 382780 338132 382844 338196
rect 386460 338132 386524 338196
rect 408172 338132 408236 338196
rect 57836 337996 57900 338060
rect 70716 337996 70780 338060
rect 60596 337860 60660 337924
rect 55996 337724 56060 337788
rect 57100 337724 57164 337788
rect 59676 337724 59740 337788
rect 63172 337724 63236 337788
rect 64276 337724 64340 337788
rect 53604 337588 53668 337652
rect 73660 337860 73724 337924
rect 78076 337860 78140 337924
rect 93348 337860 93412 337924
rect 376156 337860 376220 337924
rect 379468 337920 379532 337924
rect 379468 337864 379518 337920
rect 379518 337864 379532 337920
rect 379468 337860 379532 337864
rect 395660 337860 395724 337924
rect 398052 337860 398116 337924
rect 68324 337724 68388 337788
rect 78444 337724 78508 337788
rect 85988 337724 86052 337788
rect 88196 337724 88260 337788
rect 88748 337724 88812 337788
rect 91508 337724 91572 337788
rect 97028 337724 97092 337788
rect 103284 337724 103348 337788
rect 113404 337724 113468 337788
rect 115980 337724 116044 337788
rect 118556 337784 118620 337788
rect 118556 337728 118606 337784
rect 118606 337728 118620 337784
rect 118556 337724 118620 337728
rect 123524 337724 123588 337788
rect 125916 337724 125980 337788
rect 133460 337724 133524 337788
rect 135852 337724 135916 337788
rect 138612 337724 138676 337788
rect 143396 337784 143460 337788
rect 143396 337728 143446 337784
rect 143446 337728 143460 337784
rect 143396 337724 143460 337728
rect 145972 337724 146036 337788
rect 364196 337724 364260 337788
rect 367508 337724 367572 337788
rect 370084 337724 370148 337788
rect 373580 337724 373644 337788
rect 378548 337724 378612 337788
rect 381676 337724 381740 337788
rect 389772 337724 389836 337788
rect 392164 337724 392228 337788
rect 68692 337588 68756 337652
rect 71268 337648 71332 337652
rect 71268 337592 71318 337648
rect 71318 337592 71332 337648
rect 71268 337588 71332 337592
rect 74580 337648 74644 337652
rect 74580 337592 74630 337648
rect 74630 337592 74644 337648
rect 74580 337588 74644 337592
rect 79548 337588 79612 337652
rect 81756 337588 81820 337652
rect 83412 337588 83476 337652
rect 85252 337588 85316 337652
rect 86356 337588 86420 337652
rect 87644 337588 87708 337652
rect 89852 337588 89916 337652
rect 92244 337588 92308 337652
rect 93532 337588 93596 337652
rect 95740 337588 95804 337652
rect 97948 337588 98012 337652
rect 99236 337648 99300 337652
rect 99236 337592 99286 337648
rect 99286 337592 99300 337648
rect 99236 337588 99300 337592
rect 100892 337588 100956 337652
rect 105860 337588 105924 337652
rect 108252 337588 108316 337652
rect 111012 337588 111076 337652
rect 233188 337588 233252 337652
rect 357020 337588 357084 337652
rect 358124 337588 358188 337652
rect 359596 337588 359660 337652
rect 360516 337588 360580 337652
rect 361804 337588 361868 337652
rect 363092 337648 363156 337652
rect 363092 337592 363106 337648
rect 363106 337592 363156 337648
rect 363092 337588 363156 337592
rect 366404 337588 366468 337652
rect 368060 337588 368124 337652
rect 368980 337588 369044 337652
rect 370636 337588 370700 337652
rect 373396 337588 373460 337652
rect 374500 337588 374564 337652
rect 375788 337588 375852 337652
rect 377996 337588 378060 337652
rect 381124 337588 381188 337652
rect 385172 337588 385236 337652
rect 391060 337588 391124 337652
rect 393452 337648 393516 337652
rect 393452 337592 393466 337648
rect 393466 337592 393516 337648
rect 393452 337588 393516 337592
rect 396028 337588 396092 337652
rect 399156 337588 399220 337652
rect 401180 337588 401244 337652
rect 413324 337588 413388 337652
rect 415900 337588 415964 337652
rect 418292 337588 418356 337652
rect 420868 337648 420932 337652
rect 420868 337592 420918 337648
rect 420918 337592 420932 337648
rect 420868 337588 420932 337592
rect 428596 337588 428660 337652
rect 430988 337588 431052 337652
rect 435772 337588 435836 337652
rect 438348 337588 438412 337652
rect 445892 337588 445956 337652
rect 58204 337452 58268 337516
rect 72372 337452 72436 337516
rect 81020 337452 81084 337516
rect 82860 337452 82924 337516
rect 231900 337452 231964 337516
rect 385908 337452 385972 337516
rect 388300 337452 388364 337516
rect 356100 337316 356164 337380
rect 383516 337316 383580 337380
rect 423444 337316 423508 337380
rect 52316 337180 52380 337244
rect 61700 337180 61764 337244
rect 65380 337180 65444 337244
rect 66668 337180 66732 337244
rect 387564 337180 387628 337244
rect 410932 337180 410996 337244
rect 443316 337180 443380 337244
rect 56364 337044 56428 337108
rect 67588 337044 67652 337108
rect 141004 337044 141068 337108
rect 380572 337044 380636 337108
rect 388668 337044 388732 337108
rect 394372 337044 394436 337108
rect 433564 337044 433628 337108
rect 440924 337044 440988 337108
rect 58204 336908 58268 336972
rect 383884 336908 383948 336972
rect 393084 336908 393148 336972
rect 396580 336908 396644 336972
rect 405964 336908 406028 336972
rect 425652 336908 425716 336972
rect 70164 336772 70228 336836
rect 76052 336772 76116 336836
rect 94268 336772 94332 336836
rect 96108 336772 96172 336836
rect 120948 336772 121012 336836
rect 128492 336772 128556 336836
rect 365484 336772 365548 336836
rect 371188 336832 371252 336836
rect 371188 336776 371238 336832
rect 371238 336776 371252 336832
rect 371188 336772 371252 336776
rect 376892 336832 376956 336836
rect 376892 336776 376906 336832
rect 376906 336776 376956 336832
rect 376892 336772 376956 336776
rect 391244 336772 391308 336836
rect 398420 336772 398484 336836
rect 403572 336772 403636 336836
rect 73476 239864 73540 239868
rect 73476 239808 73490 239864
rect 73490 239808 73540 239864
rect 73476 239804 73540 239808
rect 57652 239728 57716 239732
rect 57652 239672 57702 239728
rect 57702 239672 57716 239728
rect 57652 239668 57716 239672
rect 59124 239728 59188 239732
rect 59124 239672 59174 239728
rect 59174 239672 59188 239728
rect 59124 239668 59188 239672
rect 75868 239728 75932 239732
rect 75868 239672 75882 239728
rect 75882 239672 75932 239728
rect 75868 239668 75932 239672
rect 59308 239396 59372 239460
rect 40540 47364 40604 47428
rect 40540 45460 40604 45524
rect 58204 39944 58268 39948
rect 58204 39888 58254 39944
rect 58254 39888 58268 39944
rect 58204 39884 58268 39888
rect 52316 38524 52380 38588
rect 233188 38524 233252 38588
rect 57652 38388 57716 38452
rect 231900 38388 231964 38452
rect 59124 38252 59188 38316
rect 59308 38116 59372 38180
rect 56364 37980 56428 38044
rect 53604 37844 53668 37908
rect 57836 37708 57900 37772
<< metal4 >>
rect -8726 711558 -8106 711590
rect -8726 711322 -8694 711558
rect -8458 711322 -8374 711558
rect -8138 711322 -8106 711558
rect -8726 711238 -8106 711322
rect -8726 711002 -8694 711238
rect -8458 711002 -8374 711238
rect -8138 711002 -8106 711238
rect -8726 679394 -8106 711002
rect -8726 679158 -8694 679394
rect -8458 679158 -8374 679394
rect -8138 679158 -8106 679394
rect -8726 643394 -8106 679158
rect -8726 643158 -8694 643394
rect -8458 643158 -8374 643394
rect -8138 643158 -8106 643394
rect -8726 607394 -8106 643158
rect -8726 607158 -8694 607394
rect -8458 607158 -8374 607394
rect -8138 607158 -8106 607394
rect -8726 571394 -8106 607158
rect -8726 571158 -8694 571394
rect -8458 571158 -8374 571394
rect -8138 571158 -8106 571394
rect -8726 535394 -8106 571158
rect -8726 535158 -8694 535394
rect -8458 535158 -8374 535394
rect -8138 535158 -8106 535394
rect -8726 499394 -8106 535158
rect -8726 499158 -8694 499394
rect -8458 499158 -8374 499394
rect -8138 499158 -8106 499394
rect -8726 463394 -8106 499158
rect -8726 463158 -8694 463394
rect -8458 463158 -8374 463394
rect -8138 463158 -8106 463394
rect -8726 427394 -8106 463158
rect -8726 427158 -8694 427394
rect -8458 427158 -8374 427394
rect -8138 427158 -8106 427394
rect -8726 391394 -8106 427158
rect -8726 391158 -8694 391394
rect -8458 391158 -8374 391394
rect -8138 391158 -8106 391394
rect -8726 355394 -8106 391158
rect -8726 355158 -8694 355394
rect -8458 355158 -8374 355394
rect -8138 355158 -8106 355394
rect -8726 319394 -8106 355158
rect -8726 319158 -8694 319394
rect -8458 319158 -8374 319394
rect -8138 319158 -8106 319394
rect -8726 283394 -8106 319158
rect -8726 283158 -8694 283394
rect -8458 283158 -8374 283394
rect -8138 283158 -8106 283394
rect -8726 247394 -8106 283158
rect -8726 247158 -8694 247394
rect -8458 247158 -8374 247394
rect -8138 247158 -8106 247394
rect -8726 211394 -8106 247158
rect -8726 211158 -8694 211394
rect -8458 211158 -8374 211394
rect -8138 211158 -8106 211394
rect -8726 175394 -8106 211158
rect -8726 175158 -8694 175394
rect -8458 175158 -8374 175394
rect -8138 175158 -8106 175394
rect -8726 139394 -8106 175158
rect -8726 139158 -8694 139394
rect -8458 139158 -8374 139394
rect -8138 139158 -8106 139394
rect -8726 103394 -8106 139158
rect -8726 103158 -8694 103394
rect -8458 103158 -8374 103394
rect -8138 103158 -8106 103394
rect -8726 67394 -8106 103158
rect -8726 67158 -8694 67394
rect -8458 67158 -8374 67394
rect -8138 67158 -8106 67394
rect -8726 31394 -8106 67158
rect -8726 31158 -8694 31394
rect -8458 31158 -8374 31394
rect -8138 31158 -8106 31394
rect -8726 -7066 -8106 31158
rect -7766 710598 -7146 710630
rect -7766 710362 -7734 710598
rect -7498 710362 -7414 710598
rect -7178 710362 -7146 710598
rect -7766 710278 -7146 710362
rect -7766 710042 -7734 710278
rect -7498 710042 -7414 710278
rect -7178 710042 -7146 710278
rect -7766 697394 -7146 710042
rect 11904 710598 12504 711590
rect 11904 710362 12086 710598
rect 12322 710362 12504 710598
rect 11904 710278 12504 710362
rect 11904 710042 12086 710278
rect 12322 710042 12504 710278
rect -7766 697158 -7734 697394
rect -7498 697158 -7414 697394
rect -7178 697158 -7146 697394
rect -7766 661394 -7146 697158
rect -7766 661158 -7734 661394
rect -7498 661158 -7414 661394
rect -7178 661158 -7146 661394
rect -7766 625394 -7146 661158
rect -7766 625158 -7734 625394
rect -7498 625158 -7414 625394
rect -7178 625158 -7146 625394
rect -7766 589394 -7146 625158
rect -7766 589158 -7734 589394
rect -7498 589158 -7414 589394
rect -7178 589158 -7146 589394
rect -7766 553394 -7146 589158
rect -7766 553158 -7734 553394
rect -7498 553158 -7414 553394
rect -7178 553158 -7146 553394
rect -7766 517394 -7146 553158
rect -7766 517158 -7734 517394
rect -7498 517158 -7414 517394
rect -7178 517158 -7146 517394
rect -7766 481394 -7146 517158
rect -7766 481158 -7734 481394
rect -7498 481158 -7414 481394
rect -7178 481158 -7146 481394
rect -7766 445394 -7146 481158
rect -7766 445158 -7734 445394
rect -7498 445158 -7414 445394
rect -7178 445158 -7146 445394
rect -7766 409394 -7146 445158
rect -7766 409158 -7734 409394
rect -7498 409158 -7414 409394
rect -7178 409158 -7146 409394
rect -7766 373394 -7146 409158
rect -7766 373158 -7734 373394
rect -7498 373158 -7414 373394
rect -7178 373158 -7146 373394
rect -7766 337394 -7146 373158
rect -7766 337158 -7734 337394
rect -7498 337158 -7414 337394
rect -7178 337158 -7146 337394
rect -7766 301394 -7146 337158
rect -7766 301158 -7734 301394
rect -7498 301158 -7414 301394
rect -7178 301158 -7146 301394
rect -7766 265394 -7146 301158
rect -7766 265158 -7734 265394
rect -7498 265158 -7414 265394
rect -7178 265158 -7146 265394
rect -7766 229394 -7146 265158
rect -7766 229158 -7734 229394
rect -7498 229158 -7414 229394
rect -7178 229158 -7146 229394
rect -7766 193394 -7146 229158
rect -7766 193158 -7734 193394
rect -7498 193158 -7414 193394
rect -7178 193158 -7146 193394
rect -7766 157394 -7146 193158
rect -7766 157158 -7734 157394
rect -7498 157158 -7414 157394
rect -7178 157158 -7146 157394
rect -7766 121394 -7146 157158
rect -7766 121158 -7734 121394
rect -7498 121158 -7414 121394
rect -7178 121158 -7146 121394
rect -7766 85394 -7146 121158
rect -7766 85158 -7734 85394
rect -7498 85158 -7414 85394
rect -7178 85158 -7146 85394
rect -7766 49394 -7146 85158
rect -7766 49158 -7734 49394
rect -7498 49158 -7414 49394
rect -7178 49158 -7146 49394
rect -7766 13394 -7146 49158
rect -7766 13158 -7734 13394
rect -7498 13158 -7414 13394
rect -7178 13158 -7146 13394
rect -7766 -6106 -7146 13158
rect -6806 709638 -6186 709670
rect -6806 709402 -6774 709638
rect -6538 709402 -6454 709638
rect -6218 709402 -6186 709638
rect -6806 709318 -6186 709402
rect -6806 709082 -6774 709318
rect -6538 709082 -6454 709318
rect -6218 709082 -6186 709318
rect -6806 675694 -6186 709082
rect -6806 675458 -6774 675694
rect -6538 675458 -6454 675694
rect -6218 675458 -6186 675694
rect -6806 639694 -6186 675458
rect -6806 639458 -6774 639694
rect -6538 639458 -6454 639694
rect -6218 639458 -6186 639694
rect -6806 603694 -6186 639458
rect -6806 603458 -6774 603694
rect -6538 603458 -6454 603694
rect -6218 603458 -6186 603694
rect -6806 567694 -6186 603458
rect -6806 567458 -6774 567694
rect -6538 567458 -6454 567694
rect -6218 567458 -6186 567694
rect -6806 531694 -6186 567458
rect -6806 531458 -6774 531694
rect -6538 531458 -6454 531694
rect -6218 531458 -6186 531694
rect -6806 495694 -6186 531458
rect -6806 495458 -6774 495694
rect -6538 495458 -6454 495694
rect -6218 495458 -6186 495694
rect -6806 459694 -6186 495458
rect -6806 459458 -6774 459694
rect -6538 459458 -6454 459694
rect -6218 459458 -6186 459694
rect -6806 423694 -6186 459458
rect -6806 423458 -6774 423694
rect -6538 423458 -6454 423694
rect -6218 423458 -6186 423694
rect -6806 387694 -6186 423458
rect -6806 387458 -6774 387694
rect -6538 387458 -6454 387694
rect -6218 387458 -6186 387694
rect -6806 351694 -6186 387458
rect -6806 351458 -6774 351694
rect -6538 351458 -6454 351694
rect -6218 351458 -6186 351694
rect -6806 315694 -6186 351458
rect -6806 315458 -6774 315694
rect -6538 315458 -6454 315694
rect -6218 315458 -6186 315694
rect -6806 279694 -6186 315458
rect -6806 279458 -6774 279694
rect -6538 279458 -6454 279694
rect -6218 279458 -6186 279694
rect -6806 243694 -6186 279458
rect -6806 243458 -6774 243694
rect -6538 243458 -6454 243694
rect -6218 243458 -6186 243694
rect -6806 207694 -6186 243458
rect -6806 207458 -6774 207694
rect -6538 207458 -6454 207694
rect -6218 207458 -6186 207694
rect -6806 171694 -6186 207458
rect -6806 171458 -6774 171694
rect -6538 171458 -6454 171694
rect -6218 171458 -6186 171694
rect -6806 135694 -6186 171458
rect -6806 135458 -6774 135694
rect -6538 135458 -6454 135694
rect -6218 135458 -6186 135694
rect -6806 99694 -6186 135458
rect -6806 99458 -6774 99694
rect -6538 99458 -6454 99694
rect -6218 99458 -6186 99694
rect -6806 63694 -6186 99458
rect -6806 63458 -6774 63694
rect -6538 63458 -6454 63694
rect -6218 63458 -6186 63694
rect -6806 27694 -6186 63458
rect -6806 27458 -6774 27694
rect -6538 27458 -6454 27694
rect -6218 27458 -6186 27694
rect -6806 -5146 -6186 27458
rect -5846 708678 -5226 708710
rect -5846 708442 -5814 708678
rect -5578 708442 -5494 708678
rect -5258 708442 -5226 708678
rect -5846 708358 -5226 708442
rect -5846 708122 -5814 708358
rect -5578 708122 -5494 708358
rect -5258 708122 -5226 708358
rect -5846 693694 -5226 708122
rect 8204 708678 8804 709670
rect 8204 708442 8386 708678
rect 8622 708442 8804 708678
rect 8204 708358 8804 708442
rect 8204 708122 8386 708358
rect 8622 708122 8804 708358
rect -5846 693458 -5814 693694
rect -5578 693458 -5494 693694
rect -5258 693458 -5226 693694
rect -5846 657694 -5226 693458
rect -5846 657458 -5814 657694
rect -5578 657458 -5494 657694
rect -5258 657458 -5226 657694
rect -5846 621694 -5226 657458
rect -5846 621458 -5814 621694
rect -5578 621458 -5494 621694
rect -5258 621458 -5226 621694
rect -5846 585694 -5226 621458
rect -5846 585458 -5814 585694
rect -5578 585458 -5494 585694
rect -5258 585458 -5226 585694
rect -5846 549694 -5226 585458
rect -5846 549458 -5814 549694
rect -5578 549458 -5494 549694
rect -5258 549458 -5226 549694
rect -5846 513694 -5226 549458
rect -5846 513458 -5814 513694
rect -5578 513458 -5494 513694
rect -5258 513458 -5226 513694
rect -5846 477694 -5226 513458
rect -5846 477458 -5814 477694
rect -5578 477458 -5494 477694
rect -5258 477458 -5226 477694
rect -5846 441694 -5226 477458
rect -5846 441458 -5814 441694
rect -5578 441458 -5494 441694
rect -5258 441458 -5226 441694
rect -5846 405694 -5226 441458
rect -5846 405458 -5814 405694
rect -5578 405458 -5494 405694
rect -5258 405458 -5226 405694
rect -5846 369694 -5226 405458
rect -5846 369458 -5814 369694
rect -5578 369458 -5494 369694
rect -5258 369458 -5226 369694
rect -5846 333694 -5226 369458
rect -5846 333458 -5814 333694
rect -5578 333458 -5494 333694
rect -5258 333458 -5226 333694
rect -5846 297694 -5226 333458
rect -5846 297458 -5814 297694
rect -5578 297458 -5494 297694
rect -5258 297458 -5226 297694
rect -5846 261694 -5226 297458
rect -5846 261458 -5814 261694
rect -5578 261458 -5494 261694
rect -5258 261458 -5226 261694
rect -5846 225694 -5226 261458
rect -5846 225458 -5814 225694
rect -5578 225458 -5494 225694
rect -5258 225458 -5226 225694
rect -5846 189694 -5226 225458
rect -5846 189458 -5814 189694
rect -5578 189458 -5494 189694
rect -5258 189458 -5226 189694
rect -5846 153694 -5226 189458
rect -5846 153458 -5814 153694
rect -5578 153458 -5494 153694
rect -5258 153458 -5226 153694
rect -5846 117694 -5226 153458
rect -5846 117458 -5814 117694
rect -5578 117458 -5494 117694
rect -5258 117458 -5226 117694
rect -5846 81694 -5226 117458
rect -5846 81458 -5814 81694
rect -5578 81458 -5494 81694
rect -5258 81458 -5226 81694
rect -5846 45694 -5226 81458
rect -5846 45458 -5814 45694
rect -5578 45458 -5494 45694
rect -5258 45458 -5226 45694
rect -5846 9694 -5226 45458
rect -5846 9458 -5814 9694
rect -5578 9458 -5494 9694
rect -5258 9458 -5226 9694
rect -5846 -4186 -5226 9458
rect -4886 707718 -4266 707750
rect -4886 707482 -4854 707718
rect -4618 707482 -4534 707718
rect -4298 707482 -4266 707718
rect -4886 707398 -4266 707482
rect -4886 707162 -4854 707398
rect -4618 707162 -4534 707398
rect -4298 707162 -4266 707398
rect -4886 671994 -4266 707162
rect -4886 671758 -4854 671994
rect -4618 671758 -4534 671994
rect -4298 671758 -4266 671994
rect -4886 635994 -4266 671758
rect -4886 635758 -4854 635994
rect -4618 635758 -4534 635994
rect -4298 635758 -4266 635994
rect -4886 599994 -4266 635758
rect -4886 599758 -4854 599994
rect -4618 599758 -4534 599994
rect -4298 599758 -4266 599994
rect -4886 563994 -4266 599758
rect -4886 563758 -4854 563994
rect -4618 563758 -4534 563994
rect -4298 563758 -4266 563994
rect -4886 527994 -4266 563758
rect -4886 527758 -4854 527994
rect -4618 527758 -4534 527994
rect -4298 527758 -4266 527994
rect -4886 491994 -4266 527758
rect -4886 491758 -4854 491994
rect -4618 491758 -4534 491994
rect -4298 491758 -4266 491994
rect -4886 455994 -4266 491758
rect -4886 455758 -4854 455994
rect -4618 455758 -4534 455994
rect -4298 455758 -4266 455994
rect -4886 419994 -4266 455758
rect -4886 419758 -4854 419994
rect -4618 419758 -4534 419994
rect -4298 419758 -4266 419994
rect -4886 383994 -4266 419758
rect -4886 383758 -4854 383994
rect -4618 383758 -4534 383994
rect -4298 383758 -4266 383994
rect -4886 347994 -4266 383758
rect -4886 347758 -4854 347994
rect -4618 347758 -4534 347994
rect -4298 347758 -4266 347994
rect -4886 311994 -4266 347758
rect -4886 311758 -4854 311994
rect -4618 311758 -4534 311994
rect -4298 311758 -4266 311994
rect -4886 275994 -4266 311758
rect -4886 275758 -4854 275994
rect -4618 275758 -4534 275994
rect -4298 275758 -4266 275994
rect -4886 239994 -4266 275758
rect -4886 239758 -4854 239994
rect -4618 239758 -4534 239994
rect -4298 239758 -4266 239994
rect -4886 203994 -4266 239758
rect -4886 203758 -4854 203994
rect -4618 203758 -4534 203994
rect -4298 203758 -4266 203994
rect -4886 167994 -4266 203758
rect -4886 167758 -4854 167994
rect -4618 167758 -4534 167994
rect -4298 167758 -4266 167994
rect -4886 131994 -4266 167758
rect -4886 131758 -4854 131994
rect -4618 131758 -4534 131994
rect -4298 131758 -4266 131994
rect -4886 95994 -4266 131758
rect -4886 95758 -4854 95994
rect -4618 95758 -4534 95994
rect -4298 95758 -4266 95994
rect -4886 59994 -4266 95758
rect -4886 59758 -4854 59994
rect -4618 59758 -4534 59994
rect -4298 59758 -4266 59994
rect -4886 23994 -4266 59758
rect -4886 23758 -4854 23994
rect -4618 23758 -4534 23994
rect -4298 23758 -4266 23994
rect -4886 -3226 -4266 23758
rect -3926 706758 -3306 706790
rect -3926 706522 -3894 706758
rect -3658 706522 -3574 706758
rect -3338 706522 -3306 706758
rect -3926 706438 -3306 706522
rect -3926 706202 -3894 706438
rect -3658 706202 -3574 706438
rect -3338 706202 -3306 706438
rect -3926 689994 -3306 706202
rect 4504 706758 5104 707750
rect 4504 706522 4686 706758
rect 4922 706522 5104 706758
rect 4504 706438 5104 706522
rect 4504 706202 4686 706438
rect 4922 706202 5104 706438
rect -3926 689758 -3894 689994
rect -3658 689758 -3574 689994
rect -3338 689758 -3306 689994
rect -3926 653994 -3306 689758
rect -3926 653758 -3894 653994
rect -3658 653758 -3574 653994
rect -3338 653758 -3306 653994
rect -3926 617994 -3306 653758
rect -3926 617758 -3894 617994
rect -3658 617758 -3574 617994
rect -3338 617758 -3306 617994
rect -3926 581994 -3306 617758
rect -3926 581758 -3894 581994
rect -3658 581758 -3574 581994
rect -3338 581758 -3306 581994
rect -3926 545994 -3306 581758
rect -3926 545758 -3894 545994
rect -3658 545758 -3574 545994
rect -3338 545758 -3306 545994
rect -3926 509994 -3306 545758
rect -3926 509758 -3894 509994
rect -3658 509758 -3574 509994
rect -3338 509758 -3306 509994
rect -3926 473994 -3306 509758
rect -3926 473758 -3894 473994
rect -3658 473758 -3574 473994
rect -3338 473758 -3306 473994
rect -3926 437994 -3306 473758
rect -3926 437758 -3894 437994
rect -3658 437758 -3574 437994
rect -3338 437758 -3306 437994
rect -3926 401994 -3306 437758
rect -3926 401758 -3894 401994
rect -3658 401758 -3574 401994
rect -3338 401758 -3306 401994
rect -3926 365994 -3306 401758
rect -3926 365758 -3894 365994
rect -3658 365758 -3574 365994
rect -3338 365758 -3306 365994
rect -3926 329994 -3306 365758
rect -3926 329758 -3894 329994
rect -3658 329758 -3574 329994
rect -3338 329758 -3306 329994
rect -3926 293994 -3306 329758
rect -3926 293758 -3894 293994
rect -3658 293758 -3574 293994
rect -3338 293758 -3306 293994
rect -3926 257994 -3306 293758
rect -3926 257758 -3894 257994
rect -3658 257758 -3574 257994
rect -3338 257758 -3306 257994
rect -3926 221994 -3306 257758
rect -3926 221758 -3894 221994
rect -3658 221758 -3574 221994
rect -3338 221758 -3306 221994
rect -3926 185994 -3306 221758
rect -3926 185758 -3894 185994
rect -3658 185758 -3574 185994
rect -3338 185758 -3306 185994
rect -3926 149994 -3306 185758
rect -3926 149758 -3894 149994
rect -3658 149758 -3574 149994
rect -3338 149758 -3306 149994
rect -3926 113994 -3306 149758
rect -3926 113758 -3894 113994
rect -3658 113758 -3574 113994
rect -3338 113758 -3306 113994
rect -3926 77994 -3306 113758
rect -3926 77758 -3894 77994
rect -3658 77758 -3574 77994
rect -3338 77758 -3306 77994
rect -3926 41994 -3306 77758
rect -3926 41758 -3894 41994
rect -3658 41758 -3574 41994
rect -3338 41758 -3306 41994
rect -3926 5994 -3306 41758
rect -3926 5758 -3894 5994
rect -3658 5758 -3574 5994
rect -3338 5758 -3306 5994
rect -3926 -2266 -3306 5758
rect -2966 705798 -2346 705830
rect -2966 705562 -2934 705798
rect -2698 705562 -2614 705798
rect -2378 705562 -2346 705798
rect -2966 705478 -2346 705562
rect -2966 705242 -2934 705478
rect -2698 705242 -2614 705478
rect -2378 705242 -2346 705478
rect -2966 668294 -2346 705242
rect -2966 668058 -2934 668294
rect -2698 668058 -2614 668294
rect -2378 668058 -2346 668294
rect -2966 632294 -2346 668058
rect -2966 632058 -2934 632294
rect -2698 632058 -2614 632294
rect -2378 632058 -2346 632294
rect -2966 596294 -2346 632058
rect -2966 596058 -2934 596294
rect -2698 596058 -2614 596294
rect -2378 596058 -2346 596294
rect -2966 560294 -2346 596058
rect -2966 560058 -2934 560294
rect -2698 560058 -2614 560294
rect -2378 560058 -2346 560294
rect -2966 524294 -2346 560058
rect -2966 524058 -2934 524294
rect -2698 524058 -2614 524294
rect -2378 524058 -2346 524294
rect -2966 488294 -2346 524058
rect -2966 488058 -2934 488294
rect -2698 488058 -2614 488294
rect -2378 488058 -2346 488294
rect -2966 452294 -2346 488058
rect -2966 452058 -2934 452294
rect -2698 452058 -2614 452294
rect -2378 452058 -2346 452294
rect -2966 416294 -2346 452058
rect -2966 416058 -2934 416294
rect -2698 416058 -2614 416294
rect -2378 416058 -2346 416294
rect -2966 380294 -2346 416058
rect -2966 380058 -2934 380294
rect -2698 380058 -2614 380294
rect -2378 380058 -2346 380294
rect -2966 344294 -2346 380058
rect -2966 344058 -2934 344294
rect -2698 344058 -2614 344294
rect -2378 344058 -2346 344294
rect -2966 308294 -2346 344058
rect -2966 308058 -2934 308294
rect -2698 308058 -2614 308294
rect -2378 308058 -2346 308294
rect -2966 272294 -2346 308058
rect -2966 272058 -2934 272294
rect -2698 272058 -2614 272294
rect -2378 272058 -2346 272294
rect -2966 236294 -2346 272058
rect -2966 236058 -2934 236294
rect -2698 236058 -2614 236294
rect -2378 236058 -2346 236294
rect -2966 200294 -2346 236058
rect -2966 200058 -2934 200294
rect -2698 200058 -2614 200294
rect -2378 200058 -2346 200294
rect -2966 164294 -2346 200058
rect -2966 164058 -2934 164294
rect -2698 164058 -2614 164294
rect -2378 164058 -2346 164294
rect -2966 128294 -2346 164058
rect -2966 128058 -2934 128294
rect -2698 128058 -2614 128294
rect -2378 128058 -2346 128294
rect -2966 92294 -2346 128058
rect -2966 92058 -2934 92294
rect -2698 92058 -2614 92294
rect -2378 92058 -2346 92294
rect -2966 56294 -2346 92058
rect -2966 56058 -2934 56294
rect -2698 56058 -2614 56294
rect -2378 56058 -2346 56294
rect -2966 20294 -2346 56058
rect -2966 20058 -2934 20294
rect -2698 20058 -2614 20294
rect -2378 20058 -2346 20294
rect -2966 -1306 -2346 20058
rect -2006 704838 -1386 704870
rect -2006 704602 -1974 704838
rect -1738 704602 -1654 704838
rect -1418 704602 -1386 704838
rect -2006 704518 -1386 704602
rect -2006 704282 -1974 704518
rect -1738 704282 -1654 704518
rect -1418 704282 -1386 704518
rect -2006 686294 -1386 704282
rect -2006 686058 -1974 686294
rect -1738 686058 -1654 686294
rect -1418 686058 -1386 686294
rect -2006 650294 -1386 686058
rect -2006 650058 -1974 650294
rect -1738 650058 -1654 650294
rect -1418 650058 -1386 650294
rect -2006 614294 -1386 650058
rect -2006 614058 -1974 614294
rect -1738 614058 -1654 614294
rect -1418 614058 -1386 614294
rect -2006 578294 -1386 614058
rect -2006 578058 -1974 578294
rect -1738 578058 -1654 578294
rect -1418 578058 -1386 578294
rect -2006 542294 -1386 578058
rect -2006 542058 -1974 542294
rect -1738 542058 -1654 542294
rect -1418 542058 -1386 542294
rect -2006 506294 -1386 542058
rect -2006 506058 -1974 506294
rect -1738 506058 -1654 506294
rect -1418 506058 -1386 506294
rect -2006 470294 -1386 506058
rect -2006 470058 -1974 470294
rect -1738 470058 -1654 470294
rect -1418 470058 -1386 470294
rect -2006 434294 -1386 470058
rect -2006 434058 -1974 434294
rect -1738 434058 -1654 434294
rect -1418 434058 -1386 434294
rect -2006 398294 -1386 434058
rect -2006 398058 -1974 398294
rect -1738 398058 -1654 398294
rect -1418 398058 -1386 398294
rect -2006 362294 -1386 398058
rect -2006 362058 -1974 362294
rect -1738 362058 -1654 362294
rect -1418 362058 -1386 362294
rect -2006 326294 -1386 362058
rect -2006 326058 -1974 326294
rect -1738 326058 -1654 326294
rect -1418 326058 -1386 326294
rect -2006 290294 -1386 326058
rect -2006 290058 -1974 290294
rect -1738 290058 -1654 290294
rect -1418 290058 -1386 290294
rect -2006 254294 -1386 290058
rect -2006 254058 -1974 254294
rect -1738 254058 -1654 254294
rect -1418 254058 -1386 254294
rect -2006 218294 -1386 254058
rect -2006 218058 -1974 218294
rect -1738 218058 -1654 218294
rect -1418 218058 -1386 218294
rect -2006 182294 -1386 218058
rect -2006 182058 -1974 182294
rect -1738 182058 -1654 182294
rect -1418 182058 -1386 182294
rect -2006 146294 -1386 182058
rect -2006 146058 -1974 146294
rect -1738 146058 -1654 146294
rect -1418 146058 -1386 146294
rect -2006 110294 -1386 146058
rect -2006 110058 -1974 110294
rect -1738 110058 -1654 110294
rect -1418 110058 -1386 110294
rect -2006 74294 -1386 110058
rect -2006 74058 -1974 74294
rect -1738 74058 -1654 74294
rect -1418 74058 -1386 74294
rect -2006 38294 -1386 74058
rect -2006 38058 -1974 38294
rect -1738 38058 -1654 38294
rect -1418 38058 -1386 38294
rect -2006 2294 -1386 38058
rect -2006 2058 -1974 2294
rect -1738 2058 -1654 2294
rect -1418 2058 -1386 2294
rect -2006 -346 -1386 2058
rect -2006 -582 -1974 -346
rect -1738 -582 -1654 -346
rect -1418 -582 -1386 -346
rect -2006 -666 -1386 -582
rect -2006 -902 -1974 -666
rect -1738 -902 -1654 -666
rect -1418 -902 -1386 -666
rect -2006 -934 -1386 -902
rect 804 704838 1404 705830
rect 804 704602 986 704838
rect 1222 704602 1404 704838
rect 804 704518 1404 704602
rect 804 704282 986 704518
rect 1222 704282 1404 704518
rect 804 686294 1404 704282
rect 804 686058 986 686294
rect 1222 686058 1404 686294
rect 804 650294 1404 686058
rect 804 650058 986 650294
rect 1222 650058 1404 650294
rect 804 614294 1404 650058
rect 804 614058 986 614294
rect 1222 614058 1404 614294
rect 804 578294 1404 614058
rect 804 578058 986 578294
rect 1222 578058 1404 578294
rect 804 542294 1404 578058
rect 804 542058 986 542294
rect 1222 542058 1404 542294
rect 804 506294 1404 542058
rect 804 506058 986 506294
rect 1222 506058 1404 506294
rect 804 470294 1404 506058
rect 804 470058 986 470294
rect 1222 470058 1404 470294
rect 804 434294 1404 470058
rect 804 434058 986 434294
rect 1222 434058 1404 434294
rect 804 398294 1404 434058
rect 804 398058 986 398294
rect 1222 398058 1404 398294
rect 804 362294 1404 398058
rect 804 362058 986 362294
rect 1222 362058 1404 362294
rect 804 326294 1404 362058
rect 804 326058 986 326294
rect 1222 326058 1404 326294
rect 804 290294 1404 326058
rect 804 290058 986 290294
rect 1222 290058 1404 290294
rect 804 254294 1404 290058
rect 804 254058 986 254294
rect 1222 254058 1404 254294
rect 804 218294 1404 254058
rect 804 218058 986 218294
rect 1222 218058 1404 218294
rect 804 182294 1404 218058
rect 804 182058 986 182294
rect 1222 182058 1404 182294
rect 804 146294 1404 182058
rect 804 146058 986 146294
rect 1222 146058 1404 146294
rect 804 110294 1404 146058
rect 804 110058 986 110294
rect 1222 110058 1404 110294
rect 804 74294 1404 110058
rect 804 74058 986 74294
rect 1222 74058 1404 74294
rect 804 38294 1404 74058
rect 804 38058 986 38294
rect 1222 38058 1404 38294
rect 804 2294 1404 38058
rect 804 2058 986 2294
rect 1222 2058 1404 2294
rect 804 -346 1404 2058
rect 804 -582 986 -346
rect 1222 -582 1404 -346
rect 804 -666 1404 -582
rect 804 -902 986 -666
rect 1222 -902 1404 -666
rect -2966 -1542 -2934 -1306
rect -2698 -1542 -2614 -1306
rect -2378 -1542 -2346 -1306
rect -2966 -1626 -2346 -1542
rect -2966 -1862 -2934 -1626
rect -2698 -1862 -2614 -1626
rect -2378 -1862 -2346 -1626
rect -2966 -1894 -2346 -1862
rect 804 -1894 1404 -902
rect 4504 689994 5104 706202
rect 4504 689758 4686 689994
rect 4922 689758 5104 689994
rect 4504 653994 5104 689758
rect 4504 653758 4686 653994
rect 4922 653758 5104 653994
rect 4504 617994 5104 653758
rect 4504 617758 4686 617994
rect 4922 617758 5104 617994
rect 4504 581994 5104 617758
rect 4504 581758 4686 581994
rect 4922 581758 5104 581994
rect 4504 545994 5104 581758
rect 4504 545758 4686 545994
rect 4922 545758 5104 545994
rect 4504 509994 5104 545758
rect 4504 509758 4686 509994
rect 4922 509758 5104 509994
rect 4504 473994 5104 509758
rect 4504 473758 4686 473994
rect 4922 473758 5104 473994
rect 4504 437994 5104 473758
rect 4504 437758 4686 437994
rect 4922 437758 5104 437994
rect 4504 401994 5104 437758
rect 4504 401758 4686 401994
rect 4922 401758 5104 401994
rect 4504 365994 5104 401758
rect 4504 365758 4686 365994
rect 4922 365758 5104 365994
rect 4504 329994 5104 365758
rect 4504 329758 4686 329994
rect 4922 329758 5104 329994
rect 4504 293994 5104 329758
rect 4504 293758 4686 293994
rect 4922 293758 5104 293994
rect 4504 257994 5104 293758
rect 4504 257758 4686 257994
rect 4922 257758 5104 257994
rect 4504 221994 5104 257758
rect 4504 221758 4686 221994
rect 4922 221758 5104 221994
rect 4504 185994 5104 221758
rect 4504 185758 4686 185994
rect 4922 185758 5104 185994
rect 4504 149994 5104 185758
rect 4504 149758 4686 149994
rect 4922 149758 5104 149994
rect 4504 113994 5104 149758
rect 4504 113758 4686 113994
rect 4922 113758 5104 113994
rect 4504 77994 5104 113758
rect 4504 77758 4686 77994
rect 4922 77758 5104 77994
rect 4504 41994 5104 77758
rect 4504 41758 4686 41994
rect 4922 41758 5104 41994
rect 4504 5994 5104 41758
rect 4504 5758 4686 5994
rect 4922 5758 5104 5994
rect -3926 -2502 -3894 -2266
rect -3658 -2502 -3574 -2266
rect -3338 -2502 -3306 -2266
rect -3926 -2586 -3306 -2502
rect -3926 -2822 -3894 -2586
rect -3658 -2822 -3574 -2586
rect -3338 -2822 -3306 -2586
rect -3926 -2854 -3306 -2822
rect 4504 -2266 5104 5758
rect 4504 -2502 4686 -2266
rect 4922 -2502 5104 -2266
rect 4504 -2586 5104 -2502
rect 4504 -2822 4686 -2586
rect 4922 -2822 5104 -2586
rect -4886 -3462 -4854 -3226
rect -4618 -3462 -4534 -3226
rect -4298 -3462 -4266 -3226
rect -4886 -3546 -4266 -3462
rect -4886 -3782 -4854 -3546
rect -4618 -3782 -4534 -3546
rect -4298 -3782 -4266 -3546
rect -4886 -3814 -4266 -3782
rect 4504 -3814 5104 -2822
rect 8204 693694 8804 708122
rect 8204 693458 8386 693694
rect 8622 693458 8804 693694
rect 8204 657694 8804 693458
rect 8204 657458 8386 657694
rect 8622 657458 8804 657694
rect 8204 621694 8804 657458
rect 8204 621458 8386 621694
rect 8622 621458 8804 621694
rect 8204 585694 8804 621458
rect 8204 585458 8386 585694
rect 8622 585458 8804 585694
rect 8204 549694 8804 585458
rect 8204 549458 8386 549694
rect 8622 549458 8804 549694
rect 8204 513694 8804 549458
rect 8204 513458 8386 513694
rect 8622 513458 8804 513694
rect 8204 477694 8804 513458
rect 8204 477458 8386 477694
rect 8622 477458 8804 477694
rect 8204 441694 8804 477458
rect 8204 441458 8386 441694
rect 8622 441458 8804 441694
rect 8204 405694 8804 441458
rect 8204 405458 8386 405694
rect 8622 405458 8804 405694
rect 8204 369694 8804 405458
rect 8204 369458 8386 369694
rect 8622 369458 8804 369694
rect 8204 333694 8804 369458
rect 8204 333458 8386 333694
rect 8622 333458 8804 333694
rect 8204 297694 8804 333458
rect 8204 297458 8386 297694
rect 8622 297458 8804 297694
rect 8204 261694 8804 297458
rect 8204 261458 8386 261694
rect 8622 261458 8804 261694
rect 8204 225694 8804 261458
rect 8204 225458 8386 225694
rect 8622 225458 8804 225694
rect 8204 189694 8804 225458
rect 8204 189458 8386 189694
rect 8622 189458 8804 189694
rect 8204 153694 8804 189458
rect 8204 153458 8386 153694
rect 8622 153458 8804 153694
rect 8204 117694 8804 153458
rect 8204 117458 8386 117694
rect 8622 117458 8804 117694
rect 8204 81694 8804 117458
rect 8204 81458 8386 81694
rect 8622 81458 8804 81694
rect 8204 45694 8804 81458
rect 8204 45458 8386 45694
rect 8622 45458 8804 45694
rect 8204 9694 8804 45458
rect 8204 9458 8386 9694
rect 8622 9458 8804 9694
rect -5846 -4422 -5814 -4186
rect -5578 -4422 -5494 -4186
rect -5258 -4422 -5226 -4186
rect -5846 -4506 -5226 -4422
rect -5846 -4742 -5814 -4506
rect -5578 -4742 -5494 -4506
rect -5258 -4742 -5226 -4506
rect -5846 -4774 -5226 -4742
rect 8204 -4186 8804 9458
rect 8204 -4422 8386 -4186
rect 8622 -4422 8804 -4186
rect 8204 -4506 8804 -4422
rect 8204 -4742 8386 -4506
rect 8622 -4742 8804 -4506
rect -6806 -5382 -6774 -5146
rect -6538 -5382 -6454 -5146
rect -6218 -5382 -6186 -5146
rect -6806 -5466 -6186 -5382
rect -6806 -5702 -6774 -5466
rect -6538 -5702 -6454 -5466
rect -6218 -5702 -6186 -5466
rect -6806 -5734 -6186 -5702
rect 8204 -5734 8804 -4742
rect 11904 697394 12504 710042
rect 29904 711558 30504 711590
rect 29904 711322 30086 711558
rect 30322 711322 30504 711558
rect 29904 711238 30504 711322
rect 29904 711002 30086 711238
rect 30322 711002 30504 711238
rect 26204 709638 26804 709670
rect 26204 709402 26386 709638
rect 26622 709402 26804 709638
rect 26204 709318 26804 709402
rect 26204 709082 26386 709318
rect 26622 709082 26804 709318
rect 22504 707718 23104 707750
rect 22504 707482 22686 707718
rect 22922 707482 23104 707718
rect 22504 707398 23104 707482
rect 22504 707162 22686 707398
rect 22922 707162 23104 707398
rect 11904 697158 12086 697394
rect 12322 697158 12504 697394
rect 11904 661394 12504 697158
rect 11904 661158 12086 661394
rect 12322 661158 12504 661394
rect 11904 625394 12504 661158
rect 11904 625158 12086 625394
rect 12322 625158 12504 625394
rect 11904 589394 12504 625158
rect 11904 589158 12086 589394
rect 12322 589158 12504 589394
rect 11904 553394 12504 589158
rect 11904 553158 12086 553394
rect 12322 553158 12504 553394
rect 11904 517394 12504 553158
rect 11904 517158 12086 517394
rect 12322 517158 12504 517394
rect 11904 481394 12504 517158
rect 11904 481158 12086 481394
rect 12322 481158 12504 481394
rect 11904 445394 12504 481158
rect 11904 445158 12086 445394
rect 12322 445158 12504 445394
rect 11904 409394 12504 445158
rect 11904 409158 12086 409394
rect 12322 409158 12504 409394
rect 11904 373394 12504 409158
rect 11904 373158 12086 373394
rect 12322 373158 12504 373394
rect 11904 337394 12504 373158
rect 11904 337158 12086 337394
rect 12322 337158 12504 337394
rect 11904 301394 12504 337158
rect 11904 301158 12086 301394
rect 12322 301158 12504 301394
rect 11904 265394 12504 301158
rect 11904 265158 12086 265394
rect 12322 265158 12504 265394
rect 11904 229394 12504 265158
rect 11904 229158 12086 229394
rect 12322 229158 12504 229394
rect 11904 193394 12504 229158
rect 11904 193158 12086 193394
rect 12322 193158 12504 193394
rect 11904 157394 12504 193158
rect 11904 157158 12086 157394
rect 12322 157158 12504 157394
rect 11904 121394 12504 157158
rect 11904 121158 12086 121394
rect 12322 121158 12504 121394
rect 11904 85394 12504 121158
rect 11904 85158 12086 85394
rect 12322 85158 12504 85394
rect 11904 49394 12504 85158
rect 11904 49158 12086 49394
rect 12322 49158 12504 49394
rect 11904 13394 12504 49158
rect 11904 13158 12086 13394
rect 12322 13158 12504 13394
rect -7766 -6342 -7734 -6106
rect -7498 -6342 -7414 -6106
rect -7178 -6342 -7146 -6106
rect -7766 -6426 -7146 -6342
rect -7766 -6662 -7734 -6426
rect -7498 -6662 -7414 -6426
rect -7178 -6662 -7146 -6426
rect -7766 -6694 -7146 -6662
rect 11904 -6106 12504 13158
rect 18804 705798 19404 705830
rect 18804 705562 18986 705798
rect 19222 705562 19404 705798
rect 18804 705478 19404 705562
rect 18804 705242 18986 705478
rect 19222 705242 19404 705478
rect 18804 668294 19404 705242
rect 18804 668058 18986 668294
rect 19222 668058 19404 668294
rect 18804 632294 19404 668058
rect 18804 632058 18986 632294
rect 19222 632058 19404 632294
rect 18804 596294 19404 632058
rect 18804 596058 18986 596294
rect 19222 596058 19404 596294
rect 18804 560294 19404 596058
rect 18804 560058 18986 560294
rect 19222 560058 19404 560294
rect 18804 524294 19404 560058
rect 18804 524058 18986 524294
rect 19222 524058 19404 524294
rect 18804 488294 19404 524058
rect 18804 488058 18986 488294
rect 19222 488058 19404 488294
rect 18804 452294 19404 488058
rect 18804 452058 18986 452294
rect 19222 452058 19404 452294
rect 18804 416294 19404 452058
rect 18804 416058 18986 416294
rect 19222 416058 19404 416294
rect 18804 380294 19404 416058
rect 18804 380058 18986 380294
rect 19222 380058 19404 380294
rect 18804 344294 19404 380058
rect 18804 344058 18986 344294
rect 19222 344058 19404 344294
rect 18804 308294 19404 344058
rect 18804 308058 18986 308294
rect 19222 308058 19404 308294
rect 18804 272294 19404 308058
rect 18804 272058 18986 272294
rect 19222 272058 19404 272294
rect 18804 236294 19404 272058
rect 18804 236058 18986 236294
rect 19222 236058 19404 236294
rect 18804 200294 19404 236058
rect 18804 200058 18986 200294
rect 19222 200058 19404 200294
rect 18804 164294 19404 200058
rect 18804 164058 18986 164294
rect 19222 164058 19404 164294
rect 18804 128294 19404 164058
rect 18804 128058 18986 128294
rect 19222 128058 19404 128294
rect 18804 92294 19404 128058
rect 18804 92058 18986 92294
rect 19222 92058 19404 92294
rect 18804 56294 19404 92058
rect 18804 56058 18986 56294
rect 19222 56058 19404 56294
rect 18804 20294 19404 56058
rect 18804 20058 18986 20294
rect 19222 20058 19404 20294
rect 18804 -1306 19404 20058
rect 18804 -1542 18986 -1306
rect 19222 -1542 19404 -1306
rect 18804 -1626 19404 -1542
rect 18804 -1862 18986 -1626
rect 19222 -1862 19404 -1626
rect 18804 -1894 19404 -1862
rect 22504 671994 23104 707162
rect 22504 671758 22686 671994
rect 22922 671758 23104 671994
rect 22504 635994 23104 671758
rect 22504 635758 22686 635994
rect 22922 635758 23104 635994
rect 22504 599994 23104 635758
rect 22504 599758 22686 599994
rect 22922 599758 23104 599994
rect 22504 563994 23104 599758
rect 22504 563758 22686 563994
rect 22922 563758 23104 563994
rect 22504 527994 23104 563758
rect 22504 527758 22686 527994
rect 22922 527758 23104 527994
rect 22504 491994 23104 527758
rect 22504 491758 22686 491994
rect 22922 491758 23104 491994
rect 22504 455994 23104 491758
rect 22504 455758 22686 455994
rect 22922 455758 23104 455994
rect 22504 419994 23104 455758
rect 22504 419758 22686 419994
rect 22922 419758 23104 419994
rect 22504 383994 23104 419758
rect 22504 383758 22686 383994
rect 22922 383758 23104 383994
rect 22504 347994 23104 383758
rect 22504 347758 22686 347994
rect 22922 347758 23104 347994
rect 22504 311994 23104 347758
rect 22504 311758 22686 311994
rect 22922 311758 23104 311994
rect 22504 275994 23104 311758
rect 22504 275758 22686 275994
rect 22922 275758 23104 275994
rect 22504 239994 23104 275758
rect 22504 239758 22686 239994
rect 22922 239758 23104 239994
rect 22504 203994 23104 239758
rect 22504 203758 22686 203994
rect 22922 203758 23104 203994
rect 22504 167994 23104 203758
rect 22504 167758 22686 167994
rect 22922 167758 23104 167994
rect 22504 131994 23104 167758
rect 22504 131758 22686 131994
rect 22922 131758 23104 131994
rect 22504 95994 23104 131758
rect 22504 95758 22686 95994
rect 22922 95758 23104 95994
rect 22504 59994 23104 95758
rect 22504 59758 22686 59994
rect 22922 59758 23104 59994
rect 22504 23994 23104 59758
rect 22504 23758 22686 23994
rect 22922 23758 23104 23994
rect 22504 -3226 23104 23758
rect 22504 -3462 22686 -3226
rect 22922 -3462 23104 -3226
rect 22504 -3546 23104 -3462
rect 22504 -3782 22686 -3546
rect 22922 -3782 23104 -3546
rect 22504 -3814 23104 -3782
rect 26204 675694 26804 709082
rect 26204 675458 26386 675694
rect 26622 675458 26804 675694
rect 26204 639694 26804 675458
rect 26204 639458 26386 639694
rect 26622 639458 26804 639694
rect 26204 603694 26804 639458
rect 26204 603458 26386 603694
rect 26622 603458 26804 603694
rect 26204 567694 26804 603458
rect 26204 567458 26386 567694
rect 26622 567458 26804 567694
rect 26204 531694 26804 567458
rect 26204 531458 26386 531694
rect 26622 531458 26804 531694
rect 26204 495694 26804 531458
rect 26204 495458 26386 495694
rect 26622 495458 26804 495694
rect 26204 459694 26804 495458
rect 26204 459458 26386 459694
rect 26622 459458 26804 459694
rect 26204 423694 26804 459458
rect 26204 423458 26386 423694
rect 26622 423458 26804 423694
rect 26204 387694 26804 423458
rect 26204 387458 26386 387694
rect 26622 387458 26804 387694
rect 26204 351694 26804 387458
rect 26204 351458 26386 351694
rect 26622 351458 26804 351694
rect 26204 315694 26804 351458
rect 26204 315458 26386 315694
rect 26622 315458 26804 315694
rect 26204 279694 26804 315458
rect 26204 279458 26386 279694
rect 26622 279458 26804 279694
rect 26204 243694 26804 279458
rect 26204 243458 26386 243694
rect 26622 243458 26804 243694
rect 26204 207694 26804 243458
rect 26204 207458 26386 207694
rect 26622 207458 26804 207694
rect 26204 171694 26804 207458
rect 26204 171458 26386 171694
rect 26622 171458 26804 171694
rect 26204 135694 26804 171458
rect 26204 135458 26386 135694
rect 26622 135458 26804 135694
rect 26204 99694 26804 135458
rect 26204 99458 26386 99694
rect 26622 99458 26804 99694
rect 26204 63694 26804 99458
rect 26204 63458 26386 63694
rect 26622 63458 26804 63694
rect 26204 27694 26804 63458
rect 26204 27458 26386 27694
rect 26622 27458 26804 27694
rect 26204 -5146 26804 27458
rect 26204 -5382 26386 -5146
rect 26622 -5382 26804 -5146
rect 26204 -5466 26804 -5382
rect 26204 -5702 26386 -5466
rect 26622 -5702 26804 -5466
rect 26204 -5734 26804 -5702
rect 29904 679394 30504 711002
rect 47904 710598 48504 711590
rect 47904 710362 48086 710598
rect 48322 710362 48504 710598
rect 47904 710278 48504 710362
rect 47904 710042 48086 710278
rect 48322 710042 48504 710278
rect 44204 708678 44804 709670
rect 44204 708442 44386 708678
rect 44622 708442 44804 708678
rect 44204 708358 44804 708442
rect 44204 708122 44386 708358
rect 44622 708122 44804 708358
rect 40504 706758 41104 707750
rect 40504 706522 40686 706758
rect 40922 706522 41104 706758
rect 40504 706438 41104 706522
rect 40504 706202 40686 706438
rect 40922 706202 41104 706438
rect 29904 679158 30086 679394
rect 30322 679158 30504 679394
rect 29904 643394 30504 679158
rect 29904 643158 30086 643394
rect 30322 643158 30504 643394
rect 29904 607394 30504 643158
rect 29904 607158 30086 607394
rect 30322 607158 30504 607394
rect 29904 571394 30504 607158
rect 29904 571158 30086 571394
rect 30322 571158 30504 571394
rect 29904 535394 30504 571158
rect 29904 535158 30086 535394
rect 30322 535158 30504 535394
rect 29904 499394 30504 535158
rect 29904 499158 30086 499394
rect 30322 499158 30504 499394
rect 29904 463394 30504 499158
rect 29904 463158 30086 463394
rect 30322 463158 30504 463394
rect 29904 427394 30504 463158
rect 29904 427158 30086 427394
rect 30322 427158 30504 427394
rect 29904 391394 30504 427158
rect 29904 391158 30086 391394
rect 30322 391158 30504 391394
rect 29904 355394 30504 391158
rect 29904 355158 30086 355394
rect 30322 355158 30504 355394
rect 29904 319394 30504 355158
rect 29904 319158 30086 319394
rect 30322 319158 30504 319394
rect 29904 283394 30504 319158
rect 29904 283158 30086 283394
rect 30322 283158 30504 283394
rect 29904 247394 30504 283158
rect 29904 247158 30086 247394
rect 30322 247158 30504 247394
rect 29904 211394 30504 247158
rect 29904 211158 30086 211394
rect 30322 211158 30504 211394
rect 29904 175394 30504 211158
rect 29904 175158 30086 175394
rect 30322 175158 30504 175394
rect 29904 139394 30504 175158
rect 29904 139158 30086 139394
rect 30322 139158 30504 139394
rect 29904 103394 30504 139158
rect 29904 103158 30086 103394
rect 30322 103158 30504 103394
rect 29904 67394 30504 103158
rect 29904 67158 30086 67394
rect 30322 67158 30504 67394
rect 29904 31394 30504 67158
rect 29904 31158 30086 31394
rect 30322 31158 30504 31394
rect 11904 -6342 12086 -6106
rect 12322 -6342 12504 -6106
rect 11904 -6426 12504 -6342
rect 11904 -6662 12086 -6426
rect 12322 -6662 12504 -6426
rect -8726 -7302 -8694 -7066
rect -8458 -7302 -8374 -7066
rect -8138 -7302 -8106 -7066
rect -8726 -7386 -8106 -7302
rect -8726 -7622 -8694 -7386
rect -8458 -7622 -8374 -7386
rect -8138 -7622 -8106 -7386
rect -8726 -7654 -8106 -7622
rect 11904 -7654 12504 -6662
rect 29904 -7066 30504 31158
rect 36804 704838 37404 705830
rect 36804 704602 36986 704838
rect 37222 704602 37404 704838
rect 36804 704518 37404 704602
rect 36804 704282 36986 704518
rect 37222 704282 37404 704518
rect 36804 686294 37404 704282
rect 36804 686058 36986 686294
rect 37222 686058 37404 686294
rect 36804 650294 37404 686058
rect 36804 650058 36986 650294
rect 37222 650058 37404 650294
rect 36804 614294 37404 650058
rect 36804 614058 36986 614294
rect 37222 614058 37404 614294
rect 36804 578294 37404 614058
rect 36804 578058 36986 578294
rect 37222 578058 37404 578294
rect 36804 542294 37404 578058
rect 36804 542058 36986 542294
rect 37222 542058 37404 542294
rect 36804 506294 37404 542058
rect 36804 506058 36986 506294
rect 37222 506058 37404 506294
rect 36804 470294 37404 506058
rect 36804 470058 36986 470294
rect 37222 470058 37404 470294
rect 36804 434294 37404 470058
rect 36804 434058 36986 434294
rect 37222 434058 37404 434294
rect 36804 398294 37404 434058
rect 40504 689994 41104 706202
rect 40504 689758 40686 689994
rect 40922 689758 41104 689994
rect 40504 653994 41104 689758
rect 40504 653758 40686 653994
rect 40922 653758 41104 653994
rect 40504 617994 41104 653758
rect 40504 617758 40686 617994
rect 40922 617758 41104 617994
rect 40504 581994 41104 617758
rect 40504 581758 40686 581994
rect 40922 581758 41104 581994
rect 40504 545994 41104 581758
rect 40504 545758 40686 545994
rect 40922 545758 41104 545994
rect 40504 509994 41104 545758
rect 40504 509758 40686 509994
rect 40922 509758 41104 509994
rect 40504 473994 41104 509758
rect 40504 473758 40686 473994
rect 40922 473758 41104 473994
rect 40504 437994 41104 473758
rect 40504 437758 40686 437994
rect 40922 437758 41104 437994
rect 40504 425308 41104 437758
rect 44204 693694 44804 708122
rect 44204 693458 44386 693694
rect 44622 693458 44804 693694
rect 44204 657694 44804 693458
rect 44204 657458 44386 657694
rect 44622 657458 44804 657694
rect 44204 621694 44804 657458
rect 44204 621458 44386 621694
rect 44622 621458 44804 621694
rect 44204 585694 44804 621458
rect 44204 585458 44386 585694
rect 44622 585458 44804 585694
rect 44204 549694 44804 585458
rect 44204 549458 44386 549694
rect 44622 549458 44804 549694
rect 44204 513694 44804 549458
rect 44204 513458 44386 513694
rect 44622 513458 44804 513694
rect 44204 477694 44804 513458
rect 44204 477458 44386 477694
rect 44622 477458 44804 477694
rect 44204 441694 44804 477458
rect 44204 441458 44386 441694
rect 44622 441458 44804 441694
rect 44204 425308 44804 441458
rect 47904 697394 48504 710042
rect 65904 711558 66504 711590
rect 65904 711322 66086 711558
rect 66322 711322 66504 711558
rect 65904 711238 66504 711322
rect 65904 711002 66086 711238
rect 66322 711002 66504 711238
rect 62204 709638 62804 709670
rect 62204 709402 62386 709638
rect 62622 709402 62804 709638
rect 62204 709318 62804 709402
rect 62204 709082 62386 709318
rect 62622 709082 62804 709318
rect 58504 707718 59104 707750
rect 58504 707482 58686 707718
rect 58922 707482 59104 707718
rect 58504 707398 59104 707482
rect 58504 707162 58686 707398
rect 58922 707162 59104 707398
rect 47904 697158 48086 697394
rect 48322 697158 48504 697394
rect 47904 661394 48504 697158
rect 47904 661158 48086 661394
rect 48322 661158 48504 661394
rect 47904 625394 48504 661158
rect 47904 625158 48086 625394
rect 48322 625158 48504 625394
rect 47904 589394 48504 625158
rect 47904 589158 48086 589394
rect 48322 589158 48504 589394
rect 47904 553394 48504 589158
rect 47904 553158 48086 553394
rect 48322 553158 48504 553394
rect 47904 517394 48504 553158
rect 47904 517158 48086 517394
rect 48322 517158 48504 517394
rect 47904 481394 48504 517158
rect 47904 481158 48086 481394
rect 48322 481158 48504 481394
rect 47904 445394 48504 481158
rect 47904 445158 48086 445394
rect 48322 445158 48504 445394
rect 47904 425308 48504 445158
rect 54804 705798 55404 705830
rect 54804 705562 54986 705798
rect 55222 705562 55404 705798
rect 54804 705478 55404 705562
rect 54804 705242 54986 705478
rect 55222 705242 55404 705478
rect 54804 668294 55404 705242
rect 54804 668058 54986 668294
rect 55222 668058 55404 668294
rect 54804 632294 55404 668058
rect 54804 632058 54986 632294
rect 55222 632058 55404 632294
rect 54804 596294 55404 632058
rect 54804 596058 54986 596294
rect 55222 596058 55404 596294
rect 54804 560294 55404 596058
rect 54804 560058 54986 560294
rect 55222 560058 55404 560294
rect 54804 524294 55404 560058
rect 54804 524058 54986 524294
rect 55222 524058 55404 524294
rect 54804 488294 55404 524058
rect 54804 488058 54986 488294
rect 55222 488058 55404 488294
rect 54804 452294 55404 488058
rect 54804 452058 54986 452294
rect 55222 452058 55404 452294
rect 54804 425308 55404 452058
rect 58504 671994 59104 707162
rect 58504 671758 58686 671994
rect 58922 671758 59104 671994
rect 58504 635994 59104 671758
rect 58504 635758 58686 635994
rect 58922 635758 59104 635994
rect 58504 599994 59104 635758
rect 58504 599758 58686 599994
rect 58922 599758 59104 599994
rect 58504 563994 59104 599758
rect 58504 563758 58686 563994
rect 58922 563758 59104 563994
rect 58504 527994 59104 563758
rect 58504 527758 58686 527994
rect 58922 527758 59104 527994
rect 58504 491994 59104 527758
rect 58504 491758 58686 491994
rect 58922 491758 59104 491994
rect 58504 455994 59104 491758
rect 58504 455758 58686 455994
rect 58922 455758 59104 455994
rect 58504 425308 59104 455758
rect 62204 675694 62804 709082
rect 62204 675458 62386 675694
rect 62622 675458 62804 675694
rect 62204 639694 62804 675458
rect 62204 639458 62386 639694
rect 62622 639458 62804 639694
rect 62204 603694 62804 639458
rect 62204 603458 62386 603694
rect 62622 603458 62804 603694
rect 62204 567694 62804 603458
rect 62204 567458 62386 567694
rect 62622 567458 62804 567694
rect 62204 531694 62804 567458
rect 62204 531458 62386 531694
rect 62622 531458 62804 531694
rect 62204 495694 62804 531458
rect 62204 495458 62386 495694
rect 62622 495458 62804 495694
rect 62204 459694 62804 495458
rect 62204 459458 62386 459694
rect 62622 459458 62804 459694
rect 62204 425308 62804 459458
rect 65904 679394 66504 711002
rect 83904 710598 84504 711590
rect 83904 710362 84086 710598
rect 84322 710362 84504 710598
rect 83904 710278 84504 710362
rect 83904 710042 84086 710278
rect 84322 710042 84504 710278
rect 80204 708678 80804 709670
rect 80204 708442 80386 708678
rect 80622 708442 80804 708678
rect 80204 708358 80804 708442
rect 80204 708122 80386 708358
rect 80622 708122 80804 708358
rect 76504 706758 77104 707750
rect 76504 706522 76686 706758
rect 76922 706522 77104 706758
rect 76504 706438 77104 706522
rect 76504 706202 76686 706438
rect 76922 706202 77104 706438
rect 65904 679158 66086 679394
rect 66322 679158 66504 679394
rect 65904 643394 66504 679158
rect 65904 643158 66086 643394
rect 66322 643158 66504 643394
rect 65904 607394 66504 643158
rect 65904 607158 66086 607394
rect 66322 607158 66504 607394
rect 65904 571394 66504 607158
rect 65904 571158 66086 571394
rect 66322 571158 66504 571394
rect 65904 535394 66504 571158
rect 65904 535158 66086 535394
rect 66322 535158 66504 535394
rect 65904 499394 66504 535158
rect 65904 499158 66086 499394
rect 66322 499158 66504 499394
rect 65904 463394 66504 499158
rect 65904 463158 66086 463394
rect 66322 463158 66504 463394
rect 65904 427394 66504 463158
rect 65904 427158 66086 427394
rect 66322 427158 66504 427394
rect 65904 425308 66504 427158
rect 72804 704838 73404 705830
rect 72804 704602 72986 704838
rect 73222 704602 73404 704838
rect 72804 704518 73404 704602
rect 72804 704282 72986 704518
rect 73222 704282 73404 704518
rect 72804 686294 73404 704282
rect 72804 686058 72986 686294
rect 73222 686058 73404 686294
rect 72804 650294 73404 686058
rect 72804 650058 72986 650294
rect 73222 650058 73404 650294
rect 72804 614294 73404 650058
rect 72804 614058 72986 614294
rect 73222 614058 73404 614294
rect 72804 578294 73404 614058
rect 72804 578058 72986 578294
rect 73222 578058 73404 578294
rect 72804 542294 73404 578058
rect 72804 542058 72986 542294
rect 73222 542058 73404 542294
rect 72804 506294 73404 542058
rect 72804 506058 72986 506294
rect 73222 506058 73404 506294
rect 72804 470294 73404 506058
rect 72804 470058 72986 470294
rect 73222 470058 73404 470294
rect 72804 434294 73404 470058
rect 72804 434058 72986 434294
rect 73222 434058 73404 434294
rect 72804 425308 73404 434058
rect 76504 689994 77104 706202
rect 76504 689758 76686 689994
rect 76922 689758 77104 689994
rect 76504 653994 77104 689758
rect 76504 653758 76686 653994
rect 76922 653758 77104 653994
rect 76504 617994 77104 653758
rect 76504 617758 76686 617994
rect 76922 617758 77104 617994
rect 76504 581994 77104 617758
rect 76504 581758 76686 581994
rect 76922 581758 77104 581994
rect 76504 545994 77104 581758
rect 76504 545758 76686 545994
rect 76922 545758 77104 545994
rect 76504 509994 77104 545758
rect 76504 509758 76686 509994
rect 76922 509758 77104 509994
rect 76504 473994 77104 509758
rect 76504 473758 76686 473994
rect 76922 473758 77104 473994
rect 76504 437994 77104 473758
rect 76504 437758 76686 437994
rect 76922 437758 77104 437994
rect 76504 425308 77104 437758
rect 80204 693694 80804 708122
rect 80204 693458 80386 693694
rect 80622 693458 80804 693694
rect 80204 657694 80804 693458
rect 80204 657458 80386 657694
rect 80622 657458 80804 657694
rect 80204 621694 80804 657458
rect 80204 621458 80386 621694
rect 80622 621458 80804 621694
rect 80204 585694 80804 621458
rect 80204 585458 80386 585694
rect 80622 585458 80804 585694
rect 80204 549694 80804 585458
rect 80204 549458 80386 549694
rect 80622 549458 80804 549694
rect 80204 513694 80804 549458
rect 80204 513458 80386 513694
rect 80622 513458 80804 513694
rect 80204 477694 80804 513458
rect 80204 477458 80386 477694
rect 80622 477458 80804 477694
rect 80204 441694 80804 477458
rect 80204 441458 80386 441694
rect 80622 441458 80804 441694
rect 80204 425308 80804 441458
rect 83904 697394 84504 710042
rect 101904 711558 102504 711590
rect 101904 711322 102086 711558
rect 102322 711322 102504 711558
rect 101904 711238 102504 711322
rect 101904 711002 102086 711238
rect 102322 711002 102504 711238
rect 98204 709638 98804 709670
rect 98204 709402 98386 709638
rect 98622 709402 98804 709638
rect 98204 709318 98804 709402
rect 98204 709082 98386 709318
rect 98622 709082 98804 709318
rect 94504 707718 95104 707750
rect 94504 707482 94686 707718
rect 94922 707482 95104 707718
rect 94504 707398 95104 707482
rect 94504 707162 94686 707398
rect 94922 707162 95104 707398
rect 83904 697158 84086 697394
rect 84322 697158 84504 697394
rect 83904 661394 84504 697158
rect 83904 661158 84086 661394
rect 84322 661158 84504 661394
rect 83904 625394 84504 661158
rect 83904 625158 84086 625394
rect 84322 625158 84504 625394
rect 83904 589394 84504 625158
rect 83904 589158 84086 589394
rect 84322 589158 84504 589394
rect 83904 553394 84504 589158
rect 83904 553158 84086 553394
rect 84322 553158 84504 553394
rect 83904 517394 84504 553158
rect 83904 517158 84086 517394
rect 84322 517158 84504 517394
rect 83904 481394 84504 517158
rect 83904 481158 84086 481394
rect 84322 481158 84504 481394
rect 83904 445394 84504 481158
rect 83904 445158 84086 445394
rect 84322 445158 84504 445394
rect 83904 425308 84504 445158
rect 90804 705798 91404 705830
rect 90804 705562 90986 705798
rect 91222 705562 91404 705798
rect 90804 705478 91404 705562
rect 90804 705242 90986 705478
rect 91222 705242 91404 705478
rect 90804 668294 91404 705242
rect 90804 668058 90986 668294
rect 91222 668058 91404 668294
rect 90804 632294 91404 668058
rect 90804 632058 90986 632294
rect 91222 632058 91404 632294
rect 90804 596294 91404 632058
rect 90804 596058 90986 596294
rect 91222 596058 91404 596294
rect 90804 560294 91404 596058
rect 90804 560058 90986 560294
rect 91222 560058 91404 560294
rect 90804 524294 91404 560058
rect 90804 524058 90986 524294
rect 91222 524058 91404 524294
rect 90804 488294 91404 524058
rect 90804 488058 90986 488294
rect 91222 488058 91404 488294
rect 90804 452294 91404 488058
rect 90804 452058 90986 452294
rect 91222 452058 91404 452294
rect 90804 425308 91404 452058
rect 94504 671994 95104 707162
rect 94504 671758 94686 671994
rect 94922 671758 95104 671994
rect 94504 635994 95104 671758
rect 94504 635758 94686 635994
rect 94922 635758 95104 635994
rect 94504 599994 95104 635758
rect 94504 599758 94686 599994
rect 94922 599758 95104 599994
rect 94504 563994 95104 599758
rect 94504 563758 94686 563994
rect 94922 563758 95104 563994
rect 94504 527994 95104 563758
rect 94504 527758 94686 527994
rect 94922 527758 95104 527994
rect 94504 491994 95104 527758
rect 94504 491758 94686 491994
rect 94922 491758 95104 491994
rect 94504 455994 95104 491758
rect 94504 455758 94686 455994
rect 94922 455758 95104 455994
rect 94504 425308 95104 455758
rect 98204 675694 98804 709082
rect 98204 675458 98386 675694
rect 98622 675458 98804 675694
rect 98204 639694 98804 675458
rect 98204 639458 98386 639694
rect 98622 639458 98804 639694
rect 98204 603694 98804 639458
rect 98204 603458 98386 603694
rect 98622 603458 98804 603694
rect 98204 567694 98804 603458
rect 98204 567458 98386 567694
rect 98622 567458 98804 567694
rect 98204 531694 98804 567458
rect 98204 531458 98386 531694
rect 98622 531458 98804 531694
rect 98204 495694 98804 531458
rect 98204 495458 98386 495694
rect 98622 495458 98804 495694
rect 98204 459694 98804 495458
rect 98204 459458 98386 459694
rect 98622 459458 98804 459694
rect 98204 425308 98804 459458
rect 101904 679394 102504 711002
rect 119904 710598 120504 711590
rect 119904 710362 120086 710598
rect 120322 710362 120504 710598
rect 119904 710278 120504 710362
rect 119904 710042 120086 710278
rect 120322 710042 120504 710278
rect 116204 708678 116804 709670
rect 116204 708442 116386 708678
rect 116622 708442 116804 708678
rect 116204 708358 116804 708442
rect 116204 708122 116386 708358
rect 116622 708122 116804 708358
rect 112504 706758 113104 707750
rect 112504 706522 112686 706758
rect 112922 706522 113104 706758
rect 112504 706438 113104 706522
rect 112504 706202 112686 706438
rect 112922 706202 113104 706438
rect 101904 679158 102086 679394
rect 102322 679158 102504 679394
rect 101904 643394 102504 679158
rect 101904 643158 102086 643394
rect 102322 643158 102504 643394
rect 101904 607394 102504 643158
rect 101904 607158 102086 607394
rect 102322 607158 102504 607394
rect 101904 571394 102504 607158
rect 101904 571158 102086 571394
rect 102322 571158 102504 571394
rect 101904 535394 102504 571158
rect 101904 535158 102086 535394
rect 102322 535158 102504 535394
rect 101904 499394 102504 535158
rect 101904 499158 102086 499394
rect 102322 499158 102504 499394
rect 101904 463394 102504 499158
rect 101904 463158 102086 463394
rect 102322 463158 102504 463394
rect 101904 427394 102504 463158
rect 101904 427158 102086 427394
rect 102322 427158 102504 427394
rect 101904 425308 102504 427158
rect 108804 704838 109404 705830
rect 108804 704602 108986 704838
rect 109222 704602 109404 704838
rect 108804 704518 109404 704602
rect 108804 704282 108986 704518
rect 109222 704282 109404 704518
rect 108804 686294 109404 704282
rect 108804 686058 108986 686294
rect 109222 686058 109404 686294
rect 108804 650294 109404 686058
rect 108804 650058 108986 650294
rect 109222 650058 109404 650294
rect 108804 614294 109404 650058
rect 108804 614058 108986 614294
rect 109222 614058 109404 614294
rect 108804 578294 109404 614058
rect 108804 578058 108986 578294
rect 109222 578058 109404 578294
rect 108804 542294 109404 578058
rect 108804 542058 108986 542294
rect 109222 542058 109404 542294
rect 108804 506294 109404 542058
rect 108804 506058 108986 506294
rect 109222 506058 109404 506294
rect 108804 470294 109404 506058
rect 108804 470058 108986 470294
rect 109222 470058 109404 470294
rect 108804 434294 109404 470058
rect 108804 434058 108986 434294
rect 109222 434058 109404 434294
rect 108804 425308 109404 434058
rect 112504 689994 113104 706202
rect 112504 689758 112686 689994
rect 112922 689758 113104 689994
rect 112504 653994 113104 689758
rect 112504 653758 112686 653994
rect 112922 653758 113104 653994
rect 112504 617994 113104 653758
rect 112504 617758 112686 617994
rect 112922 617758 113104 617994
rect 112504 581994 113104 617758
rect 112504 581758 112686 581994
rect 112922 581758 113104 581994
rect 112504 545994 113104 581758
rect 112504 545758 112686 545994
rect 112922 545758 113104 545994
rect 112504 509994 113104 545758
rect 112504 509758 112686 509994
rect 112922 509758 113104 509994
rect 112504 473994 113104 509758
rect 112504 473758 112686 473994
rect 112922 473758 113104 473994
rect 112504 437994 113104 473758
rect 112504 437758 112686 437994
rect 112922 437758 113104 437994
rect 112504 425308 113104 437758
rect 116204 693694 116804 708122
rect 116204 693458 116386 693694
rect 116622 693458 116804 693694
rect 116204 657694 116804 693458
rect 116204 657458 116386 657694
rect 116622 657458 116804 657694
rect 116204 621694 116804 657458
rect 116204 621458 116386 621694
rect 116622 621458 116804 621694
rect 116204 585694 116804 621458
rect 116204 585458 116386 585694
rect 116622 585458 116804 585694
rect 116204 549694 116804 585458
rect 116204 549458 116386 549694
rect 116622 549458 116804 549694
rect 116204 513694 116804 549458
rect 116204 513458 116386 513694
rect 116622 513458 116804 513694
rect 116204 477694 116804 513458
rect 116204 477458 116386 477694
rect 116622 477458 116804 477694
rect 116204 441694 116804 477458
rect 116204 441458 116386 441694
rect 116622 441458 116804 441694
rect 116204 425308 116804 441458
rect 119904 697394 120504 710042
rect 137904 711558 138504 711590
rect 137904 711322 138086 711558
rect 138322 711322 138504 711558
rect 137904 711238 138504 711322
rect 137904 711002 138086 711238
rect 138322 711002 138504 711238
rect 134204 709638 134804 709670
rect 134204 709402 134386 709638
rect 134622 709402 134804 709638
rect 134204 709318 134804 709402
rect 134204 709082 134386 709318
rect 134622 709082 134804 709318
rect 130504 707718 131104 707750
rect 130504 707482 130686 707718
rect 130922 707482 131104 707718
rect 130504 707398 131104 707482
rect 130504 707162 130686 707398
rect 130922 707162 131104 707398
rect 119904 697158 120086 697394
rect 120322 697158 120504 697394
rect 119904 661394 120504 697158
rect 119904 661158 120086 661394
rect 120322 661158 120504 661394
rect 119904 625394 120504 661158
rect 119904 625158 120086 625394
rect 120322 625158 120504 625394
rect 119904 589394 120504 625158
rect 119904 589158 120086 589394
rect 120322 589158 120504 589394
rect 119904 553394 120504 589158
rect 119904 553158 120086 553394
rect 120322 553158 120504 553394
rect 119904 517394 120504 553158
rect 119904 517158 120086 517394
rect 120322 517158 120504 517394
rect 119904 481394 120504 517158
rect 119904 481158 120086 481394
rect 120322 481158 120504 481394
rect 119904 445394 120504 481158
rect 119904 445158 120086 445394
rect 120322 445158 120504 445394
rect 119904 425308 120504 445158
rect 126804 705798 127404 705830
rect 126804 705562 126986 705798
rect 127222 705562 127404 705798
rect 126804 705478 127404 705562
rect 126804 705242 126986 705478
rect 127222 705242 127404 705478
rect 126804 668294 127404 705242
rect 126804 668058 126986 668294
rect 127222 668058 127404 668294
rect 126804 632294 127404 668058
rect 126804 632058 126986 632294
rect 127222 632058 127404 632294
rect 126804 596294 127404 632058
rect 126804 596058 126986 596294
rect 127222 596058 127404 596294
rect 126804 560294 127404 596058
rect 126804 560058 126986 560294
rect 127222 560058 127404 560294
rect 126804 524294 127404 560058
rect 126804 524058 126986 524294
rect 127222 524058 127404 524294
rect 126804 488294 127404 524058
rect 126804 488058 126986 488294
rect 127222 488058 127404 488294
rect 126804 452294 127404 488058
rect 126804 452058 126986 452294
rect 127222 452058 127404 452294
rect 126804 425308 127404 452058
rect 130504 671994 131104 707162
rect 130504 671758 130686 671994
rect 130922 671758 131104 671994
rect 130504 635994 131104 671758
rect 130504 635758 130686 635994
rect 130922 635758 131104 635994
rect 130504 599994 131104 635758
rect 130504 599758 130686 599994
rect 130922 599758 131104 599994
rect 130504 563994 131104 599758
rect 130504 563758 130686 563994
rect 130922 563758 131104 563994
rect 130504 527994 131104 563758
rect 130504 527758 130686 527994
rect 130922 527758 131104 527994
rect 130504 491994 131104 527758
rect 130504 491758 130686 491994
rect 130922 491758 131104 491994
rect 130504 455994 131104 491758
rect 130504 455758 130686 455994
rect 130922 455758 131104 455994
rect 130504 425308 131104 455758
rect 134204 675694 134804 709082
rect 134204 675458 134386 675694
rect 134622 675458 134804 675694
rect 134204 639694 134804 675458
rect 134204 639458 134386 639694
rect 134622 639458 134804 639694
rect 134204 603694 134804 639458
rect 134204 603458 134386 603694
rect 134622 603458 134804 603694
rect 134204 567694 134804 603458
rect 134204 567458 134386 567694
rect 134622 567458 134804 567694
rect 134204 531694 134804 567458
rect 134204 531458 134386 531694
rect 134622 531458 134804 531694
rect 134204 495694 134804 531458
rect 134204 495458 134386 495694
rect 134622 495458 134804 495694
rect 134204 459694 134804 495458
rect 134204 459458 134386 459694
rect 134622 459458 134804 459694
rect 134204 425308 134804 459458
rect 137904 679394 138504 711002
rect 155904 710598 156504 711590
rect 155904 710362 156086 710598
rect 156322 710362 156504 710598
rect 155904 710278 156504 710362
rect 155904 710042 156086 710278
rect 156322 710042 156504 710278
rect 152204 708678 152804 709670
rect 152204 708442 152386 708678
rect 152622 708442 152804 708678
rect 152204 708358 152804 708442
rect 152204 708122 152386 708358
rect 152622 708122 152804 708358
rect 148504 706758 149104 707750
rect 148504 706522 148686 706758
rect 148922 706522 149104 706758
rect 148504 706438 149104 706522
rect 148504 706202 148686 706438
rect 148922 706202 149104 706438
rect 137904 679158 138086 679394
rect 138322 679158 138504 679394
rect 137904 643394 138504 679158
rect 137904 643158 138086 643394
rect 138322 643158 138504 643394
rect 137904 607394 138504 643158
rect 137904 607158 138086 607394
rect 138322 607158 138504 607394
rect 137904 571394 138504 607158
rect 137904 571158 138086 571394
rect 138322 571158 138504 571394
rect 137904 535394 138504 571158
rect 137904 535158 138086 535394
rect 138322 535158 138504 535394
rect 137904 499394 138504 535158
rect 137904 499158 138086 499394
rect 138322 499158 138504 499394
rect 137904 463394 138504 499158
rect 137904 463158 138086 463394
rect 138322 463158 138504 463394
rect 137904 427394 138504 463158
rect 137904 427158 138086 427394
rect 138322 427158 138504 427394
rect 137904 425308 138504 427158
rect 144804 704838 145404 705830
rect 144804 704602 144986 704838
rect 145222 704602 145404 704838
rect 144804 704518 145404 704602
rect 144804 704282 144986 704518
rect 145222 704282 145404 704518
rect 144804 686294 145404 704282
rect 144804 686058 144986 686294
rect 145222 686058 145404 686294
rect 144804 650294 145404 686058
rect 144804 650058 144986 650294
rect 145222 650058 145404 650294
rect 144804 614294 145404 650058
rect 144804 614058 144986 614294
rect 145222 614058 145404 614294
rect 144804 578294 145404 614058
rect 144804 578058 144986 578294
rect 145222 578058 145404 578294
rect 144804 542294 145404 578058
rect 144804 542058 144986 542294
rect 145222 542058 145404 542294
rect 144804 506294 145404 542058
rect 144804 506058 144986 506294
rect 145222 506058 145404 506294
rect 144804 470294 145404 506058
rect 144804 470058 144986 470294
rect 145222 470058 145404 470294
rect 144804 434294 145404 470058
rect 144804 434058 144986 434294
rect 145222 434058 145404 434294
rect 144804 425308 145404 434058
rect 148504 689994 149104 706202
rect 148504 689758 148686 689994
rect 148922 689758 149104 689994
rect 148504 653994 149104 689758
rect 148504 653758 148686 653994
rect 148922 653758 149104 653994
rect 148504 617994 149104 653758
rect 148504 617758 148686 617994
rect 148922 617758 149104 617994
rect 148504 581994 149104 617758
rect 148504 581758 148686 581994
rect 148922 581758 149104 581994
rect 148504 545994 149104 581758
rect 148504 545758 148686 545994
rect 148922 545758 149104 545994
rect 148504 509994 149104 545758
rect 148504 509758 148686 509994
rect 148922 509758 149104 509994
rect 148504 473994 149104 509758
rect 148504 473758 148686 473994
rect 148922 473758 149104 473994
rect 148504 437994 149104 473758
rect 148504 437758 148686 437994
rect 148922 437758 149104 437994
rect 148504 425308 149104 437758
rect 152204 693694 152804 708122
rect 152204 693458 152386 693694
rect 152622 693458 152804 693694
rect 152204 657694 152804 693458
rect 152204 657458 152386 657694
rect 152622 657458 152804 657694
rect 152204 621694 152804 657458
rect 152204 621458 152386 621694
rect 152622 621458 152804 621694
rect 152204 585694 152804 621458
rect 152204 585458 152386 585694
rect 152622 585458 152804 585694
rect 152204 549694 152804 585458
rect 152204 549458 152386 549694
rect 152622 549458 152804 549694
rect 152204 513694 152804 549458
rect 152204 513458 152386 513694
rect 152622 513458 152804 513694
rect 152204 477694 152804 513458
rect 152204 477458 152386 477694
rect 152622 477458 152804 477694
rect 152204 441694 152804 477458
rect 152204 441458 152386 441694
rect 152622 441458 152804 441694
rect 152204 425308 152804 441458
rect 155904 697394 156504 710042
rect 173904 711558 174504 711590
rect 173904 711322 174086 711558
rect 174322 711322 174504 711558
rect 173904 711238 174504 711322
rect 173904 711002 174086 711238
rect 174322 711002 174504 711238
rect 170204 709638 170804 709670
rect 170204 709402 170386 709638
rect 170622 709402 170804 709638
rect 170204 709318 170804 709402
rect 170204 709082 170386 709318
rect 170622 709082 170804 709318
rect 166504 707718 167104 707750
rect 166504 707482 166686 707718
rect 166922 707482 167104 707718
rect 166504 707398 167104 707482
rect 166504 707162 166686 707398
rect 166922 707162 167104 707398
rect 155904 697158 156086 697394
rect 156322 697158 156504 697394
rect 155904 661394 156504 697158
rect 155904 661158 156086 661394
rect 156322 661158 156504 661394
rect 155904 625394 156504 661158
rect 155904 625158 156086 625394
rect 156322 625158 156504 625394
rect 155904 589394 156504 625158
rect 155904 589158 156086 589394
rect 156322 589158 156504 589394
rect 155904 553394 156504 589158
rect 155904 553158 156086 553394
rect 156322 553158 156504 553394
rect 155904 517394 156504 553158
rect 155904 517158 156086 517394
rect 156322 517158 156504 517394
rect 155904 481394 156504 517158
rect 155904 481158 156086 481394
rect 156322 481158 156504 481394
rect 155904 445394 156504 481158
rect 155904 445158 156086 445394
rect 156322 445158 156504 445394
rect 155904 425308 156504 445158
rect 162804 705798 163404 705830
rect 162804 705562 162986 705798
rect 163222 705562 163404 705798
rect 162804 705478 163404 705562
rect 162804 705242 162986 705478
rect 163222 705242 163404 705478
rect 162804 668294 163404 705242
rect 162804 668058 162986 668294
rect 163222 668058 163404 668294
rect 162804 632294 163404 668058
rect 162804 632058 162986 632294
rect 163222 632058 163404 632294
rect 162804 596294 163404 632058
rect 162804 596058 162986 596294
rect 163222 596058 163404 596294
rect 162804 560294 163404 596058
rect 162804 560058 162986 560294
rect 163222 560058 163404 560294
rect 162804 524294 163404 560058
rect 162804 524058 162986 524294
rect 163222 524058 163404 524294
rect 162804 488294 163404 524058
rect 162804 488058 162986 488294
rect 163222 488058 163404 488294
rect 162804 452294 163404 488058
rect 162804 452058 162986 452294
rect 163222 452058 163404 452294
rect 162804 425308 163404 452058
rect 166504 671994 167104 707162
rect 166504 671758 166686 671994
rect 166922 671758 167104 671994
rect 166504 635994 167104 671758
rect 166504 635758 166686 635994
rect 166922 635758 167104 635994
rect 166504 599994 167104 635758
rect 166504 599758 166686 599994
rect 166922 599758 167104 599994
rect 166504 563994 167104 599758
rect 166504 563758 166686 563994
rect 166922 563758 167104 563994
rect 166504 527994 167104 563758
rect 166504 527758 166686 527994
rect 166922 527758 167104 527994
rect 166504 491994 167104 527758
rect 166504 491758 166686 491994
rect 166922 491758 167104 491994
rect 166504 455994 167104 491758
rect 166504 455758 166686 455994
rect 166922 455758 167104 455994
rect 166504 425308 167104 455758
rect 170204 675694 170804 709082
rect 170204 675458 170386 675694
rect 170622 675458 170804 675694
rect 170204 639694 170804 675458
rect 170204 639458 170386 639694
rect 170622 639458 170804 639694
rect 170204 603694 170804 639458
rect 170204 603458 170386 603694
rect 170622 603458 170804 603694
rect 170204 567694 170804 603458
rect 170204 567458 170386 567694
rect 170622 567458 170804 567694
rect 170204 531694 170804 567458
rect 170204 531458 170386 531694
rect 170622 531458 170804 531694
rect 170204 495694 170804 531458
rect 170204 495458 170386 495694
rect 170622 495458 170804 495694
rect 170204 459694 170804 495458
rect 170204 459458 170386 459694
rect 170622 459458 170804 459694
rect 170204 425308 170804 459458
rect 173904 679394 174504 711002
rect 191904 710598 192504 711590
rect 191904 710362 192086 710598
rect 192322 710362 192504 710598
rect 191904 710278 192504 710362
rect 191904 710042 192086 710278
rect 192322 710042 192504 710278
rect 188204 708678 188804 709670
rect 188204 708442 188386 708678
rect 188622 708442 188804 708678
rect 188204 708358 188804 708442
rect 188204 708122 188386 708358
rect 188622 708122 188804 708358
rect 184504 706758 185104 707750
rect 184504 706522 184686 706758
rect 184922 706522 185104 706758
rect 184504 706438 185104 706522
rect 184504 706202 184686 706438
rect 184922 706202 185104 706438
rect 173904 679158 174086 679394
rect 174322 679158 174504 679394
rect 173904 643394 174504 679158
rect 173904 643158 174086 643394
rect 174322 643158 174504 643394
rect 173904 607394 174504 643158
rect 173904 607158 174086 607394
rect 174322 607158 174504 607394
rect 173904 571394 174504 607158
rect 173904 571158 174086 571394
rect 174322 571158 174504 571394
rect 173904 535394 174504 571158
rect 173904 535158 174086 535394
rect 174322 535158 174504 535394
rect 173904 499394 174504 535158
rect 173904 499158 174086 499394
rect 174322 499158 174504 499394
rect 173904 463394 174504 499158
rect 173904 463158 174086 463394
rect 174322 463158 174504 463394
rect 173904 427394 174504 463158
rect 173904 427158 174086 427394
rect 174322 427158 174504 427394
rect 173904 425308 174504 427158
rect 180804 704838 181404 705830
rect 180804 704602 180986 704838
rect 181222 704602 181404 704838
rect 180804 704518 181404 704602
rect 180804 704282 180986 704518
rect 181222 704282 181404 704518
rect 180804 686294 181404 704282
rect 180804 686058 180986 686294
rect 181222 686058 181404 686294
rect 180804 650294 181404 686058
rect 180804 650058 180986 650294
rect 181222 650058 181404 650294
rect 180804 614294 181404 650058
rect 180804 614058 180986 614294
rect 181222 614058 181404 614294
rect 180804 578294 181404 614058
rect 180804 578058 180986 578294
rect 181222 578058 181404 578294
rect 180804 542294 181404 578058
rect 180804 542058 180986 542294
rect 181222 542058 181404 542294
rect 180804 506294 181404 542058
rect 180804 506058 180986 506294
rect 181222 506058 181404 506294
rect 180804 470294 181404 506058
rect 180804 470058 180986 470294
rect 181222 470058 181404 470294
rect 180804 434294 181404 470058
rect 180804 434058 180986 434294
rect 181222 434058 181404 434294
rect 40272 416294 40620 416476
rect 40272 416058 40328 416294
rect 40564 416058 40620 416294
rect 40272 415876 40620 416058
rect 176000 416294 176348 416476
rect 176000 416058 176056 416294
rect 176292 416058 176348 416294
rect 176000 415876 176348 416058
rect 36804 398058 36986 398294
rect 37222 398058 37404 398294
rect 36804 362294 37404 398058
rect 40952 398294 41300 398476
rect 40952 398058 41008 398294
rect 41244 398058 41300 398294
rect 40952 397876 41300 398058
rect 175320 398294 175668 398476
rect 175320 398058 175376 398294
rect 175612 398058 175668 398294
rect 175320 397876 175668 398058
rect 180804 398294 181404 434058
rect 180804 398058 180986 398294
rect 181222 398058 181404 398294
rect 40272 380294 40620 380476
rect 40272 380058 40328 380294
rect 40564 380058 40620 380294
rect 40272 379876 40620 380058
rect 176000 380294 176348 380476
rect 176000 380058 176056 380294
rect 176292 380058 176348 380294
rect 176000 379876 176348 380058
rect 36804 362058 36986 362294
rect 37222 362058 37404 362294
rect 36804 326294 37404 362058
rect 40952 362294 41300 362476
rect 40952 362058 41008 362294
rect 41244 362058 41300 362294
rect 40952 361876 41300 362058
rect 175320 362294 175668 362476
rect 175320 362058 175376 362294
rect 175612 362058 175668 362294
rect 175320 361876 175668 362058
rect 180804 362294 181404 398058
rect 180804 362058 180986 362294
rect 181222 362058 181404 362294
rect 40272 344294 40620 344476
rect 40272 344058 40328 344294
rect 40564 344058 40620 344294
rect 40272 343876 40620 344058
rect 176000 344294 176348 344476
rect 176000 344058 176056 344294
rect 176292 344058 176348 344294
rect 176000 343876 176348 344058
rect 93534 340076 93622 340136
rect 56056 339690 56116 340000
rect 57144 339690 57204 340000
rect 58232 339690 58292 340000
rect 55998 339630 56116 339690
rect 57102 339630 57204 339690
rect 58206 339630 58292 339690
rect 59592 339690 59652 340000
rect 60544 339690 60604 340000
rect 61768 339690 61828 340000
rect 59592 339630 59738 339690
rect 60544 339630 60658 339690
rect 36804 326058 36986 326294
rect 37222 326058 37404 326294
rect 36804 290294 37404 326058
rect 36804 290058 36986 290294
rect 37222 290058 37404 290294
rect 36804 254294 37404 290058
rect 36804 254058 36986 254294
rect 37222 254058 37404 254294
rect 36804 218294 37404 254058
rect 40504 329994 41104 338000
rect 40504 329758 40686 329994
rect 40922 329758 41104 329994
rect 40504 293994 41104 329758
rect 40504 293758 40686 293994
rect 40922 293758 41104 293994
rect 40504 257994 41104 293758
rect 40504 257758 40686 257994
rect 40922 257758 41104 257994
rect 40504 242304 41104 257758
rect 44204 333694 44804 338000
rect 44204 333458 44386 333694
rect 44622 333458 44804 333694
rect 44204 297694 44804 333458
rect 44204 297458 44386 297694
rect 44622 297458 44804 297694
rect 44204 261694 44804 297458
rect 44204 261458 44386 261694
rect 44622 261458 44804 261694
rect 44204 242304 44804 261458
rect 47904 337394 48504 338000
rect 53603 337652 53669 337653
rect 53603 337588 53604 337652
rect 53668 337588 53669 337652
rect 53603 337587 53669 337588
rect 47904 337158 48086 337394
rect 48322 337158 48504 337394
rect 52315 337244 52381 337245
rect 52315 337180 52316 337244
rect 52380 337180 52381 337244
rect 52315 337179 52381 337180
rect 47904 301394 48504 337158
rect 47904 301158 48086 301394
rect 48322 301158 48504 301394
rect 47904 265394 48504 301158
rect 47904 265158 48086 265394
rect 48322 265158 48504 265394
rect 47904 242304 48504 265158
rect 36804 218058 36986 218294
rect 37222 218058 37404 218294
rect 36804 182294 37404 218058
rect 44208 218294 44528 218476
rect 44208 218058 44250 218294
rect 44486 218058 44528 218294
rect 44208 217876 44528 218058
rect 36804 182058 36986 182294
rect 37222 182058 37404 182294
rect 36804 146294 37404 182058
rect 44208 182294 44528 182476
rect 44208 182058 44250 182294
rect 44486 182058 44528 182294
rect 44208 181876 44528 182058
rect 36804 146058 36986 146294
rect 37222 146058 37404 146294
rect 36804 110294 37404 146058
rect 44208 146294 44528 146476
rect 44208 146058 44250 146294
rect 44486 146058 44528 146294
rect 44208 145876 44528 146058
rect 36804 110058 36986 110294
rect 37222 110058 37404 110294
rect 36804 74294 37404 110058
rect 44208 110294 44528 110476
rect 44208 110058 44250 110294
rect 44486 110058 44528 110294
rect 44208 109876 44528 110058
rect 36804 74058 36986 74294
rect 37222 74058 37404 74294
rect 36804 38294 37404 74058
rect 44208 74294 44528 74476
rect 44208 74058 44250 74294
rect 44486 74058 44528 74294
rect 44208 73876 44528 74058
rect 40539 47428 40605 47429
rect 40539 47364 40540 47428
rect 40604 47364 40605 47428
rect 40539 47363 40605 47364
rect 40542 45525 40602 47363
rect 40539 45524 40605 45525
rect 40539 45460 40540 45524
rect 40604 45460 40605 45524
rect 40539 45459 40605 45460
rect 52318 38589 52378 337179
rect 52315 38588 52381 38589
rect 52315 38524 52316 38588
rect 52380 38524 52381 38588
rect 52315 38523 52381 38524
rect 36804 38058 36986 38294
rect 37222 38058 37404 38294
rect 36804 2294 37404 38058
rect 36804 2058 36986 2294
rect 37222 2058 37404 2294
rect 36804 -346 37404 2058
rect 36804 -582 36986 -346
rect 37222 -582 37404 -346
rect 36804 -666 37404 -582
rect 36804 -902 36986 -666
rect 37222 -902 37404 -666
rect 36804 -1894 37404 -902
rect 40504 5994 41104 38000
rect 40504 5758 40686 5994
rect 40922 5758 41104 5994
rect 40504 -2266 41104 5758
rect 40504 -2502 40686 -2266
rect 40922 -2502 41104 -2266
rect 40504 -2586 41104 -2502
rect 40504 -2822 40686 -2586
rect 40922 -2822 41104 -2586
rect 40504 -3814 41104 -2822
rect 44204 9694 44804 38000
rect 44204 9458 44386 9694
rect 44622 9458 44804 9694
rect 44204 -4186 44804 9458
rect 44204 -4422 44386 -4186
rect 44622 -4422 44804 -4186
rect 44204 -4506 44804 -4422
rect 44204 -4742 44386 -4506
rect 44622 -4742 44804 -4506
rect 44204 -5734 44804 -4742
rect 47904 13394 48504 38000
rect 53606 37909 53666 337587
rect 54804 308294 55404 338000
rect 55998 337789 56058 339630
rect 57102 337789 57162 339630
rect 57835 338060 57901 338061
rect 57835 337996 57836 338060
rect 57900 337996 57901 338060
rect 57835 337995 57901 337996
rect 55995 337788 56061 337789
rect 55995 337724 55996 337788
rect 56060 337724 56061 337788
rect 55995 337723 56061 337724
rect 57099 337788 57165 337789
rect 57099 337724 57100 337788
rect 57164 337724 57165 337788
rect 57099 337723 57165 337724
rect 56363 337108 56429 337109
rect 56363 337044 56364 337108
rect 56428 337044 56429 337108
rect 56363 337043 56429 337044
rect 54804 308058 54986 308294
rect 55222 308058 55404 308294
rect 54804 272294 55404 308058
rect 54804 272058 54986 272294
rect 55222 272058 55404 272294
rect 54804 242304 55404 272058
rect 56366 38045 56426 337043
rect 57651 239732 57717 239733
rect 57651 239668 57652 239732
rect 57716 239668 57717 239732
rect 57651 239667 57717 239668
rect 57654 38453 57714 239667
rect 57651 38452 57717 38453
rect 57651 38388 57652 38452
rect 57716 38388 57717 38452
rect 57651 38387 57717 38388
rect 56363 38044 56429 38045
rect 53603 37908 53669 37909
rect 53603 37844 53604 37908
rect 53668 37844 53669 37908
rect 53603 37843 53669 37844
rect 47904 13158 48086 13394
rect 48322 13158 48504 13394
rect 29904 -7302 30086 -7066
rect 30322 -7302 30504 -7066
rect 29904 -7386 30504 -7302
rect 29904 -7622 30086 -7386
rect 30322 -7622 30504 -7386
rect 29904 -7654 30504 -7622
rect 47904 -6106 48504 13158
rect 54804 20294 55404 38000
rect 56363 37980 56364 38044
rect 56428 37980 56429 38044
rect 56363 37979 56429 37980
rect 57838 37773 57898 337995
rect 58206 337517 58266 339630
rect 58203 337516 58269 337517
rect 58203 337452 58204 337516
rect 58268 337452 58269 337516
rect 58203 337451 58269 337452
rect 58203 336972 58269 336973
rect 58203 336908 58204 336972
rect 58268 336908 58269 336972
rect 58203 336907 58269 336908
rect 58206 39949 58266 336907
rect 58504 311994 59104 338000
rect 59678 337789 59738 339630
rect 60598 337925 60658 339630
rect 61702 339630 61828 339690
rect 63128 339690 63188 340000
rect 64216 339690 64276 340000
rect 65440 339690 65500 340000
rect 63128 339630 63234 339690
rect 64216 339630 64338 339690
rect 60595 337924 60661 337925
rect 60595 337860 60596 337924
rect 60660 337860 60661 337924
rect 60595 337859 60661 337860
rect 59675 337788 59741 337789
rect 59675 337724 59676 337788
rect 59740 337724 59741 337788
rect 59675 337723 59741 337724
rect 61702 337245 61762 339630
rect 61699 337244 61765 337245
rect 61699 337180 61700 337244
rect 61764 337180 61765 337244
rect 61699 337179 61765 337180
rect 58504 311758 58686 311994
rect 58922 311758 59104 311994
rect 58504 275994 59104 311758
rect 58504 275758 58686 275994
rect 58922 275758 59104 275994
rect 58504 242304 59104 275758
rect 62204 315694 62804 338000
rect 63174 337789 63234 339630
rect 64278 337789 64338 339630
rect 65382 339630 65500 339690
rect 66528 339690 66588 340000
rect 67616 339690 67676 340000
rect 66528 339630 66730 339690
rect 63171 337788 63237 337789
rect 63171 337724 63172 337788
rect 63236 337724 63237 337788
rect 63171 337723 63237 337724
rect 64275 337788 64341 337789
rect 64275 337724 64276 337788
rect 64340 337724 64341 337788
rect 64275 337723 64341 337724
rect 65382 337245 65442 339630
rect 65379 337244 65445 337245
rect 65379 337180 65380 337244
rect 65444 337180 65445 337244
rect 65379 337179 65445 337180
rect 62204 315458 62386 315694
rect 62622 315458 62804 315694
rect 62204 279694 62804 315458
rect 62204 279458 62386 279694
rect 62622 279458 62804 279694
rect 62204 243694 62804 279458
rect 62204 243458 62386 243694
rect 62622 243458 62804 243694
rect 62204 242304 62804 243458
rect 65904 319394 66504 338000
rect 66670 337245 66730 339630
rect 67590 339630 67676 339690
rect 68296 339690 68356 340000
rect 68704 339690 68764 340000
rect 68296 339630 68386 339690
rect 66667 337244 66733 337245
rect 66667 337180 66668 337244
rect 66732 337180 66733 337244
rect 66667 337179 66733 337180
rect 67590 337109 67650 339630
rect 68326 337789 68386 339630
rect 68694 339630 68764 339690
rect 70064 339690 70124 340000
rect 70744 339690 70804 340000
rect 71288 339690 71348 340000
rect 72376 339690 72436 340000
rect 70064 339630 70226 339690
rect 68323 337788 68389 337789
rect 68323 337724 68324 337788
rect 68388 337724 68389 337788
rect 68323 337723 68389 337724
rect 68694 337653 68754 339630
rect 68691 337652 68757 337653
rect 68691 337588 68692 337652
rect 68756 337588 68757 337652
rect 68691 337587 68757 337588
rect 67587 337108 67653 337109
rect 67587 337044 67588 337108
rect 67652 337044 67653 337108
rect 67587 337043 67653 337044
rect 70166 336837 70226 339630
rect 70718 339630 70804 339690
rect 71270 339630 71348 339690
rect 72374 339630 72436 339690
rect 73464 339690 73524 340000
rect 73600 339690 73660 340000
rect 74552 339690 74612 340000
rect 75912 339690 75972 340000
rect 73464 339630 73538 339690
rect 73600 339630 73722 339690
rect 74552 339630 74642 339690
rect 70718 338061 70778 339630
rect 70715 338060 70781 338061
rect 70715 337996 70716 338060
rect 70780 337996 70781 338060
rect 70715 337995 70781 337996
rect 71270 337653 71330 339630
rect 71267 337652 71333 337653
rect 71267 337588 71268 337652
rect 71332 337588 71333 337652
rect 71267 337587 71333 337588
rect 72374 337517 72434 339630
rect 72371 337516 72437 337517
rect 72371 337452 72372 337516
rect 72436 337452 72437 337516
rect 72371 337451 72437 337452
rect 70163 336836 70229 336837
rect 70163 336772 70164 336836
rect 70228 336772 70229 336836
rect 70163 336771 70229 336772
rect 65904 319158 66086 319394
rect 66322 319158 66504 319394
rect 65904 283394 66504 319158
rect 65904 283158 66086 283394
rect 66322 283158 66504 283394
rect 65904 247394 66504 283158
rect 65904 247158 66086 247394
rect 66322 247158 66504 247394
rect 65904 242304 66504 247158
rect 72804 326294 73404 338000
rect 72804 326058 72986 326294
rect 73222 326058 73404 326294
rect 72804 290294 73404 326058
rect 72804 290058 72986 290294
rect 73222 290058 73404 290294
rect 72804 254294 73404 290058
rect 72804 254058 72986 254294
rect 73222 254058 73404 254294
rect 72804 242304 73404 254058
rect 73478 239869 73538 339630
rect 73662 337925 73722 339630
rect 73659 337924 73725 337925
rect 73659 337860 73660 337924
rect 73724 337860 73725 337924
rect 73659 337859 73725 337860
rect 74582 337653 74642 339630
rect 75870 339630 75972 339690
rect 76048 339690 76108 340000
rect 77000 339690 77060 340000
rect 78088 339690 78148 340000
rect 78496 339690 78556 340000
rect 76048 339630 76114 339690
rect 74579 337652 74645 337653
rect 74579 337588 74580 337652
rect 74644 337588 74645 337652
rect 74579 337587 74645 337588
rect 73475 239868 73541 239869
rect 73475 239804 73476 239868
rect 73540 239804 73541 239868
rect 73475 239803 73541 239804
rect 75870 239733 75930 339630
rect 76054 336837 76114 339630
rect 76974 339630 77060 339690
rect 78078 339630 78148 339690
rect 78446 339630 78556 339690
rect 79448 339690 79508 340000
rect 80672 339690 80732 340000
rect 81080 339690 81140 340000
rect 81760 339690 81820 340000
rect 79448 339630 79610 339690
rect 76974 338197 77034 339630
rect 76971 338196 77037 338197
rect 76971 338132 76972 338196
rect 77036 338132 77037 338196
rect 76971 338131 77037 338132
rect 76051 336836 76117 336837
rect 76051 336772 76052 336836
rect 76116 336772 76117 336836
rect 76051 336771 76117 336772
rect 76504 329994 77104 338000
rect 78078 337925 78138 339630
rect 78075 337924 78141 337925
rect 78075 337860 78076 337924
rect 78140 337860 78141 337924
rect 78075 337859 78141 337860
rect 78446 337789 78506 339630
rect 78443 337788 78509 337789
rect 78443 337724 78444 337788
rect 78508 337724 78509 337788
rect 78443 337723 78509 337724
rect 79550 337653 79610 339630
rect 80654 339630 80732 339690
rect 81022 339630 81140 339690
rect 81758 339630 81820 339690
rect 82848 339690 82908 340000
rect 83528 339690 83588 340000
rect 82848 339630 82922 339690
rect 80654 338197 80714 339630
rect 80651 338196 80717 338197
rect 80651 338132 80652 338196
rect 80716 338132 80717 338196
rect 80651 338131 80717 338132
rect 79547 337652 79613 337653
rect 79547 337588 79548 337652
rect 79612 337588 79613 337652
rect 79547 337587 79613 337588
rect 76504 329758 76686 329994
rect 76922 329758 77104 329994
rect 76504 293994 77104 329758
rect 76504 293758 76686 293994
rect 76922 293758 77104 293994
rect 76504 257994 77104 293758
rect 76504 257758 76686 257994
rect 76922 257758 77104 257994
rect 76504 242304 77104 257758
rect 80204 333694 80804 338000
rect 81022 337517 81082 339630
rect 81758 337653 81818 339630
rect 81755 337652 81821 337653
rect 81755 337588 81756 337652
rect 81820 337588 81821 337652
rect 81755 337587 81821 337588
rect 82862 337517 82922 339630
rect 83414 339630 83588 339690
rect 83936 339690 83996 340000
rect 85296 339690 85356 340000
rect 83936 339630 84026 339690
rect 83414 337653 83474 339630
rect 83966 338197 84026 339630
rect 85254 339630 85356 339690
rect 85976 339690 86036 340000
rect 86384 339690 86444 340000
rect 85976 339630 86050 339690
rect 83963 338196 84029 338197
rect 83963 338132 83964 338196
rect 84028 338132 84029 338196
rect 83963 338131 84029 338132
rect 83411 337652 83477 337653
rect 83411 337588 83412 337652
rect 83476 337588 83477 337652
rect 83411 337587 83477 337588
rect 81019 337516 81085 337517
rect 81019 337452 81020 337516
rect 81084 337452 81085 337516
rect 81019 337451 81085 337452
rect 82859 337516 82925 337517
rect 82859 337452 82860 337516
rect 82924 337452 82925 337516
rect 82859 337451 82925 337452
rect 80204 333458 80386 333694
rect 80622 333458 80804 333694
rect 80204 297694 80804 333458
rect 80204 297458 80386 297694
rect 80622 297458 80804 297694
rect 80204 261694 80804 297458
rect 80204 261458 80386 261694
rect 80622 261458 80804 261694
rect 80204 242304 80804 261458
rect 83904 337394 84504 338000
rect 85254 337653 85314 339630
rect 85990 337789 86050 339630
rect 86358 339630 86444 339690
rect 87608 339690 87668 340000
rect 88288 339690 88348 340000
rect 87608 339630 87706 339690
rect 85987 337788 86053 337789
rect 85987 337724 85988 337788
rect 86052 337724 86053 337788
rect 85987 337723 86053 337724
rect 86358 337653 86418 339630
rect 87646 337653 87706 339630
rect 88198 339630 88348 339690
rect 88696 339690 88756 340000
rect 89784 339690 89844 340000
rect 91008 339690 91068 340000
rect 88696 339630 88810 339690
rect 89784 339630 89914 339690
rect 88198 337789 88258 339630
rect 88750 337789 88810 339630
rect 88195 337788 88261 337789
rect 88195 337724 88196 337788
rect 88260 337724 88261 337788
rect 88195 337723 88261 337724
rect 88747 337788 88813 337789
rect 88747 337724 88748 337788
rect 88812 337724 88813 337788
rect 88747 337723 88813 337724
rect 89854 337653 89914 339630
rect 90958 339630 91068 339690
rect 91144 339690 91204 340000
rect 92232 339690 92292 340000
rect 93320 339690 93380 340000
rect 91144 339630 91570 339690
rect 92232 339630 92306 339690
rect 93320 339630 93410 339690
rect 90958 338197 91018 339630
rect 90955 338196 91021 338197
rect 90955 338132 90956 338196
rect 91020 338132 91021 338196
rect 90955 338131 91021 338132
rect 85251 337652 85317 337653
rect 85251 337588 85252 337652
rect 85316 337588 85317 337652
rect 85251 337587 85317 337588
rect 86355 337652 86421 337653
rect 86355 337588 86356 337652
rect 86420 337588 86421 337652
rect 86355 337587 86421 337588
rect 87643 337652 87709 337653
rect 87643 337588 87644 337652
rect 87708 337588 87709 337652
rect 87643 337587 87709 337588
rect 89851 337652 89917 337653
rect 89851 337588 89852 337652
rect 89916 337588 89917 337652
rect 89851 337587 89917 337588
rect 83904 337158 84086 337394
rect 84322 337158 84504 337394
rect 83904 301394 84504 337158
rect 83904 301158 84086 301394
rect 84322 301158 84504 301394
rect 83904 265394 84504 301158
rect 83904 265158 84086 265394
rect 84322 265158 84504 265394
rect 83904 242304 84504 265158
rect 90804 308294 91404 338000
rect 91510 337789 91570 339630
rect 91507 337788 91573 337789
rect 91507 337724 91508 337788
rect 91572 337724 91573 337788
rect 91507 337723 91573 337724
rect 92246 337653 92306 339630
rect 93350 337925 93410 339630
rect 93347 337924 93413 337925
rect 93347 337860 93348 337924
rect 93412 337860 93413 337924
rect 93347 337859 93413 337860
rect 93534 337653 93594 340076
rect 94408 339690 94468 340000
rect 95768 339690 95828 340000
rect 94270 339630 94468 339690
rect 95742 339630 95828 339690
rect 96040 339690 96100 340000
rect 96992 339690 97052 340000
rect 98080 339690 98140 340000
rect 96040 339630 96170 339690
rect 96992 339630 97090 339690
rect 92243 337652 92309 337653
rect 92243 337588 92244 337652
rect 92308 337588 92309 337652
rect 92243 337587 92309 337588
rect 93531 337652 93597 337653
rect 93531 337588 93532 337652
rect 93596 337588 93597 337652
rect 93531 337587 93597 337588
rect 94270 336837 94330 339630
rect 94267 336836 94333 336837
rect 94267 336772 94268 336836
rect 94332 336772 94333 336836
rect 94267 336771 94333 336772
rect 90804 308058 90986 308294
rect 91222 308058 91404 308294
rect 90804 272294 91404 308058
rect 90804 272058 90986 272294
rect 91222 272058 91404 272294
rect 90804 242304 91404 272058
rect 94504 311994 95104 338000
rect 95742 337653 95802 339630
rect 95739 337652 95805 337653
rect 95739 337588 95740 337652
rect 95804 337588 95805 337652
rect 95739 337587 95805 337588
rect 96110 336837 96170 339630
rect 97030 337789 97090 339630
rect 97950 339630 98140 339690
rect 98488 339690 98548 340000
rect 99168 339690 99228 340000
rect 100936 339690 100996 340000
rect 103520 339690 103580 340000
rect 105968 339690 106028 340000
rect 108280 339690 108340 340000
rect 98488 339630 98562 339690
rect 99168 339630 99298 339690
rect 97027 337788 97093 337789
rect 97027 337724 97028 337788
rect 97092 337724 97093 337788
rect 97027 337723 97093 337724
rect 97950 337653 98010 339630
rect 98502 338197 98562 339630
rect 98499 338196 98565 338197
rect 98499 338132 98500 338196
rect 98564 338132 98565 338196
rect 98499 338131 98565 338132
rect 97947 337652 98013 337653
rect 97947 337588 97948 337652
rect 98012 337588 98013 337652
rect 97947 337587 98013 337588
rect 96107 336836 96173 336837
rect 96107 336772 96108 336836
rect 96172 336772 96173 336836
rect 96107 336771 96173 336772
rect 94504 311758 94686 311994
rect 94922 311758 95104 311994
rect 94504 275994 95104 311758
rect 94504 275758 94686 275994
rect 94922 275758 95104 275994
rect 94504 242304 95104 275758
rect 98204 315694 98804 338000
rect 99238 337653 99298 339630
rect 100894 339630 100996 339690
rect 103286 339630 103580 339690
rect 105862 339630 106028 339690
rect 108254 339630 108340 339690
rect 111000 339690 111060 340000
rect 113448 339690 113508 340000
rect 111000 339630 111074 339690
rect 100894 337653 100954 339630
rect 99235 337652 99301 337653
rect 99235 337588 99236 337652
rect 99300 337588 99301 337652
rect 99235 337587 99301 337588
rect 100891 337652 100957 337653
rect 100891 337588 100892 337652
rect 100956 337588 100957 337652
rect 100891 337587 100957 337588
rect 98204 315458 98386 315694
rect 98622 315458 98804 315694
rect 98204 279694 98804 315458
rect 98204 279458 98386 279694
rect 98622 279458 98804 279694
rect 98204 243694 98804 279458
rect 98204 243458 98386 243694
rect 98622 243458 98804 243694
rect 98204 242304 98804 243458
rect 101904 319394 102504 338000
rect 103286 337789 103346 339630
rect 103283 337788 103349 337789
rect 103283 337724 103284 337788
rect 103348 337724 103349 337788
rect 103283 337723 103349 337724
rect 105862 337653 105922 339630
rect 108254 337653 108314 339630
rect 105859 337652 105925 337653
rect 105859 337588 105860 337652
rect 105924 337588 105925 337652
rect 105859 337587 105925 337588
rect 108251 337652 108317 337653
rect 108251 337588 108252 337652
rect 108316 337588 108317 337652
rect 108251 337587 108317 337588
rect 101904 319158 102086 319394
rect 102322 319158 102504 319394
rect 101904 283394 102504 319158
rect 101904 283158 102086 283394
rect 102322 283158 102504 283394
rect 101904 247394 102504 283158
rect 101904 247158 102086 247394
rect 102322 247158 102504 247394
rect 101904 242304 102504 247158
rect 108804 326294 109404 338000
rect 111014 337653 111074 339630
rect 113406 339630 113508 339690
rect 115896 339690 115956 340000
rect 118480 339690 118540 340000
rect 120928 339690 120988 340000
rect 123512 339690 123572 340000
rect 125960 339690 126020 340000
rect 128544 339690 128604 340000
rect 115896 339630 116042 339690
rect 118480 339630 118618 339690
rect 120928 339630 121010 339690
rect 123512 339630 123586 339690
rect 111011 337652 111077 337653
rect 111011 337588 111012 337652
rect 111076 337588 111077 337652
rect 111011 337587 111077 337588
rect 108804 326058 108986 326294
rect 109222 326058 109404 326294
rect 108804 290294 109404 326058
rect 108804 290058 108986 290294
rect 109222 290058 109404 290294
rect 108804 254294 109404 290058
rect 108804 254058 108986 254294
rect 109222 254058 109404 254294
rect 108804 242304 109404 254058
rect 112504 329994 113104 338000
rect 113406 337789 113466 339630
rect 115982 337789 116042 339630
rect 113403 337788 113469 337789
rect 113403 337724 113404 337788
rect 113468 337724 113469 337788
rect 113403 337723 113469 337724
rect 115979 337788 116045 337789
rect 115979 337724 115980 337788
rect 116044 337724 116045 337788
rect 115979 337723 116045 337724
rect 112504 329758 112686 329994
rect 112922 329758 113104 329994
rect 112504 293994 113104 329758
rect 112504 293758 112686 293994
rect 112922 293758 113104 293994
rect 112504 257994 113104 293758
rect 112504 257758 112686 257994
rect 112922 257758 113104 257994
rect 112504 242304 113104 257758
rect 116204 333694 116804 338000
rect 118558 337789 118618 339630
rect 118555 337788 118621 337789
rect 118555 337724 118556 337788
rect 118620 337724 118621 337788
rect 118555 337723 118621 337724
rect 116204 333458 116386 333694
rect 116622 333458 116804 333694
rect 116204 297694 116804 333458
rect 116204 297458 116386 297694
rect 116622 297458 116804 297694
rect 116204 261694 116804 297458
rect 116204 261458 116386 261694
rect 116622 261458 116804 261694
rect 116204 242304 116804 261458
rect 119904 337394 120504 338000
rect 119904 337158 120086 337394
rect 120322 337158 120504 337394
rect 119904 301394 120504 337158
rect 120950 336837 121010 339630
rect 123526 337789 123586 339630
rect 125918 339630 126020 339690
rect 128494 339630 128604 339690
rect 130992 339690 131052 340000
rect 133440 339690 133500 340000
rect 135888 339690 135948 340000
rect 130992 339630 131130 339690
rect 133440 339630 133522 339690
rect 125918 337789 125978 339630
rect 123523 337788 123589 337789
rect 123523 337724 123524 337788
rect 123588 337724 123589 337788
rect 123523 337723 123589 337724
rect 125915 337788 125981 337789
rect 125915 337724 125916 337788
rect 125980 337724 125981 337788
rect 125915 337723 125981 337724
rect 120947 336836 121013 336837
rect 120947 336772 120948 336836
rect 121012 336772 121013 336836
rect 120947 336771 121013 336772
rect 119904 301158 120086 301394
rect 120322 301158 120504 301394
rect 119904 265394 120504 301158
rect 119904 265158 120086 265394
rect 120322 265158 120504 265394
rect 119904 242304 120504 265158
rect 126804 308294 127404 338000
rect 128494 336837 128554 339630
rect 131070 338197 131130 339630
rect 131067 338196 131133 338197
rect 131067 338132 131068 338196
rect 131132 338132 131133 338196
rect 131067 338131 131133 338132
rect 128491 336836 128557 336837
rect 128491 336772 128492 336836
rect 128556 336772 128557 336836
rect 128491 336771 128557 336772
rect 126804 308058 126986 308294
rect 127222 308058 127404 308294
rect 126804 272294 127404 308058
rect 126804 272058 126986 272294
rect 127222 272058 127404 272294
rect 126804 242304 127404 272058
rect 130504 311994 131104 338000
rect 133462 337789 133522 339630
rect 135854 339630 135948 339690
rect 138472 339690 138532 340000
rect 140920 339690 140980 340000
rect 143368 339690 143428 340000
rect 145952 339690 146012 340000
rect 138472 339630 138674 339690
rect 140920 339630 141066 339690
rect 143368 339630 143458 339690
rect 145952 339630 146034 339690
rect 133459 337788 133525 337789
rect 133459 337724 133460 337788
rect 133524 337724 133525 337788
rect 133459 337723 133525 337724
rect 130504 311758 130686 311994
rect 130922 311758 131104 311994
rect 130504 275994 131104 311758
rect 130504 275758 130686 275994
rect 130922 275758 131104 275994
rect 130504 242304 131104 275758
rect 134204 315694 134804 338000
rect 135854 337789 135914 339630
rect 135851 337788 135917 337789
rect 135851 337724 135852 337788
rect 135916 337724 135917 337788
rect 135851 337723 135917 337724
rect 134204 315458 134386 315694
rect 134622 315458 134804 315694
rect 134204 279694 134804 315458
rect 134204 279458 134386 279694
rect 134622 279458 134804 279694
rect 134204 243694 134804 279458
rect 134204 243458 134386 243694
rect 134622 243458 134804 243694
rect 134204 242304 134804 243458
rect 137904 319394 138504 338000
rect 138614 337789 138674 339630
rect 138611 337788 138677 337789
rect 138611 337724 138612 337788
rect 138676 337724 138677 337788
rect 138611 337723 138677 337724
rect 141006 337109 141066 339630
rect 143398 337789 143458 339630
rect 143395 337788 143461 337789
rect 143395 337724 143396 337788
rect 143460 337724 143461 337788
rect 143395 337723 143461 337724
rect 141003 337108 141069 337109
rect 141003 337044 141004 337108
rect 141068 337044 141069 337108
rect 141003 337043 141069 337044
rect 137904 319158 138086 319394
rect 138322 319158 138504 319394
rect 137904 283394 138504 319158
rect 137904 283158 138086 283394
rect 138322 283158 138504 283394
rect 137904 247394 138504 283158
rect 137904 247158 138086 247394
rect 138322 247158 138504 247394
rect 137904 242304 138504 247158
rect 144804 326294 145404 338000
rect 145974 337789 146034 339630
rect 145971 337788 146037 337789
rect 145971 337724 145972 337788
rect 146036 337724 146037 337788
rect 145971 337723 146037 337724
rect 144804 326058 144986 326294
rect 145222 326058 145404 326294
rect 144804 290294 145404 326058
rect 144804 290058 144986 290294
rect 145222 290058 145404 290294
rect 144804 254294 145404 290058
rect 144804 254058 144986 254294
rect 145222 254058 145404 254294
rect 144804 242304 145404 254058
rect 148504 329994 149104 338000
rect 148504 329758 148686 329994
rect 148922 329758 149104 329994
rect 148504 293994 149104 329758
rect 148504 293758 148686 293994
rect 148922 293758 149104 293994
rect 148504 257994 149104 293758
rect 148504 257758 148686 257994
rect 148922 257758 149104 257994
rect 148504 242304 149104 257758
rect 152204 333694 152804 338000
rect 152204 333458 152386 333694
rect 152622 333458 152804 333694
rect 152204 297694 152804 333458
rect 152204 297458 152386 297694
rect 152622 297458 152804 297694
rect 152204 261694 152804 297458
rect 152204 261458 152386 261694
rect 152622 261458 152804 261694
rect 152204 242304 152804 261458
rect 155904 337394 156504 338000
rect 155904 337158 156086 337394
rect 156322 337158 156504 337394
rect 155904 301394 156504 337158
rect 155904 301158 156086 301394
rect 156322 301158 156504 301394
rect 155904 265394 156504 301158
rect 155904 265158 156086 265394
rect 156322 265158 156504 265394
rect 155904 242304 156504 265158
rect 162804 308294 163404 338000
rect 162804 308058 162986 308294
rect 163222 308058 163404 308294
rect 162804 272294 163404 308058
rect 162804 272058 162986 272294
rect 163222 272058 163404 272294
rect 162804 242304 163404 272058
rect 166504 311994 167104 338000
rect 166504 311758 166686 311994
rect 166922 311758 167104 311994
rect 166504 275994 167104 311758
rect 166504 275758 166686 275994
rect 166922 275758 167104 275994
rect 166504 242304 167104 275758
rect 170204 315694 170804 338000
rect 170204 315458 170386 315694
rect 170622 315458 170804 315694
rect 170204 279694 170804 315458
rect 170204 279458 170386 279694
rect 170622 279458 170804 279694
rect 170204 243694 170804 279458
rect 170204 243458 170386 243694
rect 170622 243458 170804 243694
rect 170204 242304 170804 243458
rect 173904 319394 174504 338000
rect 173904 319158 174086 319394
rect 174322 319158 174504 319394
rect 173904 283394 174504 319158
rect 173904 283158 174086 283394
rect 174322 283158 174504 283394
rect 173904 247394 174504 283158
rect 173904 247158 174086 247394
rect 174322 247158 174504 247394
rect 173904 242304 174504 247158
rect 180804 326294 181404 362058
rect 180804 326058 180986 326294
rect 181222 326058 181404 326294
rect 180804 290294 181404 326058
rect 180804 290058 180986 290294
rect 181222 290058 181404 290294
rect 180804 254294 181404 290058
rect 180804 254058 180986 254294
rect 181222 254058 181404 254294
rect 180804 242304 181404 254058
rect 184504 689994 185104 706202
rect 184504 689758 184686 689994
rect 184922 689758 185104 689994
rect 184504 653994 185104 689758
rect 184504 653758 184686 653994
rect 184922 653758 185104 653994
rect 184504 617994 185104 653758
rect 184504 617758 184686 617994
rect 184922 617758 185104 617994
rect 184504 581994 185104 617758
rect 184504 581758 184686 581994
rect 184922 581758 185104 581994
rect 184504 545994 185104 581758
rect 184504 545758 184686 545994
rect 184922 545758 185104 545994
rect 184504 509994 185104 545758
rect 184504 509758 184686 509994
rect 184922 509758 185104 509994
rect 184504 473994 185104 509758
rect 184504 473758 184686 473994
rect 184922 473758 185104 473994
rect 184504 437994 185104 473758
rect 184504 437758 184686 437994
rect 184922 437758 185104 437994
rect 184504 401994 185104 437758
rect 184504 401758 184686 401994
rect 184922 401758 185104 401994
rect 184504 365994 185104 401758
rect 184504 365758 184686 365994
rect 184922 365758 185104 365994
rect 184504 329994 185104 365758
rect 184504 329758 184686 329994
rect 184922 329758 185104 329994
rect 184504 293994 185104 329758
rect 184504 293758 184686 293994
rect 184922 293758 185104 293994
rect 184504 257994 185104 293758
rect 184504 257758 184686 257994
rect 184922 257758 185104 257994
rect 184504 242304 185104 257758
rect 188204 693694 188804 708122
rect 188204 693458 188386 693694
rect 188622 693458 188804 693694
rect 188204 657694 188804 693458
rect 188204 657458 188386 657694
rect 188622 657458 188804 657694
rect 188204 621694 188804 657458
rect 188204 621458 188386 621694
rect 188622 621458 188804 621694
rect 188204 585694 188804 621458
rect 188204 585458 188386 585694
rect 188622 585458 188804 585694
rect 188204 549694 188804 585458
rect 188204 549458 188386 549694
rect 188622 549458 188804 549694
rect 188204 513694 188804 549458
rect 188204 513458 188386 513694
rect 188622 513458 188804 513694
rect 188204 477694 188804 513458
rect 188204 477458 188386 477694
rect 188622 477458 188804 477694
rect 188204 441694 188804 477458
rect 188204 441458 188386 441694
rect 188622 441458 188804 441694
rect 188204 405694 188804 441458
rect 188204 405458 188386 405694
rect 188622 405458 188804 405694
rect 188204 369694 188804 405458
rect 188204 369458 188386 369694
rect 188622 369458 188804 369694
rect 188204 333694 188804 369458
rect 188204 333458 188386 333694
rect 188622 333458 188804 333694
rect 188204 297694 188804 333458
rect 188204 297458 188386 297694
rect 188622 297458 188804 297694
rect 188204 261694 188804 297458
rect 188204 261458 188386 261694
rect 188622 261458 188804 261694
rect 188204 242304 188804 261458
rect 191904 697394 192504 710042
rect 209904 711558 210504 711590
rect 209904 711322 210086 711558
rect 210322 711322 210504 711558
rect 209904 711238 210504 711322
rect 209904 711002 210086 711238
rect 210322 711002 210504 711238
rect 206204 709638 206804 709670
rect 206204 709402 206386 709638
rect 206622 709402 206804 709638
rect 206204 709318 206804 709402
rect 206204 709082 206386 709318
rect 206622 709082 206804 709318
rect 202504 707718 203104 707750
rect 202504 707482 202686 707718
rect 202922 707482 203104 707718
rect 202504 707398 203104 707482
rect 202504 707162 202686 707398
rect 202922 707162 203104 707398
rect 191904 697158 192086 697394
rect 192322 697158 192504 697394
rect 191904 661394 192504 697158
rect 191904 661158 192086 661394
rect 192322 661158 192504 661394
rect 191904 625394 192504 661158
rect 191904 625158 192086 625394
rect 192322 625158 192504 625394
rect 191904 589394 192504 625158
rect 191904 589158 192086 589394
rect 192322 589158 192504 589394
rect 191904 553394 192504 589158
rect 191904 553158 192086 553394
rect 192322 553158 192504 553394
rect 191904 517394 192504 553158
rect 191904 517158 192086 517394
rect 192322 517158 192504 517394
rect 191904 481394 192504 517158
rect 191904 481158 192086 481394
rect 192322 481158 192504 481394
rect 191904 445394 192504 481158
rect 191904 445158 192086 445394
rect 192322 445158 192504 445394
rect 191904 409394 192504 445158
rect 191904 409158 192086 409394
rect 192322 409158 192504 409394
rect 191904 373394 192504 409158
rect 191904 373158 192086 373394
rect 192322 373158 192504 373394
rect 191904 337394 192504 373158
rect 191904 337158 192086 337394
rect 192322 337158 192504 337394
rect 191904 301394 192504 337158
rect 191904 301158 192086 301394
rect 192322 301158 192504 301394
rect 191904 265394 192504 301158
rect 191904 265158 192086 265394
rect 192322 265158 192504 265394
rect 191904 242304 192504 265158
rect 198804 705798 199404 705830
rect 198804 705562 198986 705798
rect 199222 705562 199404 705798
rect 198804 705478 199404 705562
rect 198804 705242 198986 705478
rect 199222 705242 199404 705478
rect 198804 668294 199404 705242
rect 198804 668058 198986 668294
rect 199222 668058 199404 668294
rect 198804 632294 199404 668058
rect 198804 632058 198986 632294
rect 199222 632058 199404 632294
rect 198804 596294 199404 632058
rect 198804 596058 198986 596294
rect 199222 596058 199404 596294
rect 198804 560294 199404 596058
rect 198804 560058 198986 560294
rect 199222 560058 199404 560294
rect 198804 524294 199404 560058
rect 198804 524058 198986 524294
rect 199222 524058 199404 524294
rect 198804 488294 199404 524058
rect 198804 488058 198986 488294
rect 199222 488058 199404 488294
rect 198804 452294 199404 488058
rect 198804 452058 198986 452294
rect 199222 452058 199404 452294
rect 198804 416294 199404 452058
rect 198804 416058 198986 416294
rect 199222 416058 199404 416294
rect 198804 380294 199404 416058
rect 198804 380058 198986 380294
rect 199222 380058 199404 380294
rect 198804 344294 199404 380058
rect 198804 344058 198986 344294
rect 199222 344058 199404 344294
rect 198804 308294 199404 344058
rect 198804 308058 198986 308294
rect 199222 308058 199404 308294
rect 198804 272294 199404 308058
rect 198804 272058 198986 272294
rect 199222 272058 199404 272294
rect 198804 242304 199404 272058
rect 202504 671994 203104 707162
rect 202504 671758 202686 671994
rect 202922 671758 203104 671994
rect 202504 635994 203104 671758
rect 202504 635758 202686 635994
rect 202922 635758 203104 635994
rect 202504 599994 203104 635758
rect 202504 599758 202686 599994
rect 202922 599758 203104 599994
rect 202504 563994 203104 599758
rect 202504 563758 202686 563994
rect 202922 563758 203104 563994
rect 202504 527994 203104 563758
rect 202504 527758 202686 527994
rect 202922 527758 203104 527994
rect 202504 491994 203104 527758
rect 202504 491758 202686 491994
rect 202922 491758 203104 491994
rect 202504 455994 203104 491758
rect 202504 455758 202686 455994
rect 202922 455758 203104 455994
rect 202504 419994 203104 455758
rect 202504 419758 202686 419994
rect 202922 419758 203104 419994
rect 202504 383994 203104 419758
rect 202504 383758 202686 383994
rect 202922 383758 203104 383994
rect 202504 347994 203104 383758
rect 202504 347758 202686 347994
rect 202922 347758 203104 347994
rect 202504 311994 203104 347758
rect 202504 311758 202686 311994
rect 202922 311758 203104 311994
rect 202504 275994 203104 311758
rect 202504 275758 202686 275994
rect 202922 275758 203104 275994
rect 202504 242304 203104 275758
rect 206204 675694 206804 709082
rect 206204 675458 206386 675694
rect 206622 675458 206804 675694
rect 206204 639694 206804 675458
rect 206204 639458 206386 639694
rect 206622 639458 206804 639694
rect 206204 603694 206804 639458
rect 206204 603458 206386 603694
rect 206622 603458 206804 603694
rect 206204 567694 206804 603458
rect 206204 567458 206386 567694
rect 206622 567458 206804 567694
rect 206204 531694 206804 567458
rect 206204 531458 206386 531694
rect 206622 531458 206804 531694
rect 206204 495694 206804 531458
rect 206204 495458 206386 495694
rect 206622 495458 206804 495694
rect 206204 459694 206804 495458
rect 206204 459458 206386 459694
rect 206622 459458 206804 459694
rect 206204 423694 206804 459458
rect 206204 423458 206386 423694
rect 206622 423458 206804 423694
rect 206204 387694 206804 423458
rect 206204 387458 206386 387694
rect 206622 387458 206804 387694
rect 206204 351694 206804 387458
rect 206204 351458 206386 351694
rect 206622 351458 206804 351694
rect 206204 315694 206804 351458
rect 206204 315458 206386 315694
rect 206622 315458 206804 315694
rect 206204 279694 206804 315458
rect 206204 279458 206386 279694
rect 206622 279458 206804 279694
rect 206204 243694 206804 279458
rect 206204 243458 206386 243694
rect 206622 243458 206804 243694
rect 206204 242304 206804 243458
rect 209904 679394 210504 711002
rect 227904 710598 228504 711590
rect 227904 710362 228086 710598
rect 228322 710362 228504 710598
rect 227904 710278 228504 710362
rect 227904 710042 228086 710278
rect 228322 710042 228504 710278
rect 224204 708678 224804 709670
rect 224204 708442 224386 708678
rect 224622 708442 224804 708678
rect 224204 708358 224804 708442
rect 224204 708122 224386 708358
rect 224622 708122 224804 708358
rect 220504 706758 221104 707750
rect 220504 706522 220686 706758
rect 220922 706522 221104 706758
rect 220504 706438 221104 706522
rect 220504 706202 220686 706438
rect 220922 706202 221104 706438
rect 209904 679158 210086 679394
rect 210322 679158 210504 679394
rect 209904 643394 210504 679158
rect 209904 643158 210086 643394
rect 210322 643158 210504 643394
rect 209904 607394 210504 643158
rect 209904 607158 210086 607394
rect 210322 607158 210504 607394
rect 209904 571394 210504 607158
rect 209904 571158 210086 571394
rect 210322 571158 210504 571394
rect 209904 535394 210504 571158
rect 209904 535158 210086 535394
rect 210322 535158 210504 535394
rect 209904 499394 210504 535158
rect 209904 499158 210086 499394
rect 210322 499158 210504 499394
rect 209904 463394 210504 499158
rect 209904 463158 210086 463394
rect 210322 463158 210504 463394
rect 209904 427394 210504 463158
rect 209904 427158 210086 427394
rect 210322 427158 210504 427394
rect 209904 391394 210504 427158
rect 209904 391158 210086 391394
rect 210322 391158 210504 391394
rect 209904 355394 210504 391158
rect 209904 355158 210086 355394
rect 210322 355158 210504 355394
rect 209904 319394 210504 355158
rect 209904 319158 210086 319394
rect 210322 319158 210504 319394
rect 209904 283394 210504 319158
rect 209904 283158 210086 283394
rect 210322 283158 210504 283394
rect 209904 247394 210504 283158
rect 209904 247158 210086 247394
rect 210322 247158 210504 247394
rect 209904 242304 210504 247158
rect 216804 704838 217404 705830
rect 216804 704602 216986 704838
rect 217222 704602 217404 704838
rect 216804 704518 217404 704602
rect 216804 704282 216986 704518
rect 217222 704282 217404 704518
rect 216804 686294 217404 704282
rect 216804 686058 216986 686294
rect 217222 686058 217404 686294
rect 216804 650294 217404 686058
rect 216804 650058 216986 650294
rect 217222 650058 217404 650294
rect 216804 614294 217404 650058
rect 216804 614058 216986 614294
rect 217222 614058 217404 614294
rect 216804 578294 217404 614058
rect 216804 578058 216986 578294
rect 217222 578058 217404 578294
rect 216804 542294 217404 578058
rect 216804 542058 216986 542294
rect 217222 542058 217404 542294
rect 216804 506294 217404 542058
rect 216804 506058 216986 506294
rect 217222 506058 217404 506294
rect 216804 470294 217404 506058
rect 216804 470058 216986 470294
rect 217222 470058 217404 470294
rect 216804 434294 217404 470058
rect 216804 434058 216986 434294
rect 217222 434058 217404 434294
rect 216804 398294 217404 434058
rect 216804 398058 216986 398294
rect 217222 398058 217404 398294
rect 216804 362294 217404 398058
rect 216804 362058 216986 362294
rect 217222 362058 217404 362294
rect 216804 326294 217404 362058
rect 216804 326058 216986 326294
rect 217222 326058 217404 326294
rect 216804 290294 217404 326058
rect 216804 290058 216986 290294
rect 217222 290058 217404 290294
rect 216804 254294 217404 290058
rect 216804 254058 216986 254294
rect 217222 254058 217404 254294
rect 216804 242304 217404 254058
rect 220504 689994 221104 706202
rect 220504 689758 220686 689994
rect 220922 689758 221104 689994
rect 220504 653994 221104 689758
rect 220504 653758 220686 653994
rect 220922 653758 221104 653994
rect 220504 617994 221104 653758
rect 220504 617758 220686 617994
rect 220922 617758 221104 617994
rect 220504 581994 221104 617758
rect 220504 581758 220686 581994
rect 220922 581758 221104 581994
rect 220504 545994 221104 581758
rect 220504 545758 220686 545994
rect 220922 545758 221104 545994
rect 220504 509994 221104 545758
rect 220504 509758 220686 509994
rect 220922 509758 221104 509994
rect 220504 473994 221104 509758
rect 220504 473758 220686 473994
rect 220922 473758 221104 473994
rect 220504 437994 221104 473758
rect 220504 437758 220686 437994
rect 220922 437758 221104 437994
rect 220504 401994 221104 437758
rect 220504 401758 220686 401994
rect 220922 401758 221104 401994
rect 220504 365994 221104 401758
rect 220504 365758 220686 365994
rect 220922 365758 221104 365994
rect 220504 329994 221104 365758
rect 220504 329758 220686 329994
rect 220922 329758 221104 329994
rect 220504 293994 221104 329758
rect 220504 293758 220686 293994
rect 220922 293758 221104 293994
rect 220504 257994 221104 293758
rect 220504 257758 220686 257994
rect 220922 257758 221104 257994
rect 220504 242304 221104 257758
rect 224204 693694 224804 708122
rect 224204 693458 224386 693694
rect 224622 693458 224804 693694
rect 224204 657694 224804 693458
rect 224204 657458 224386 657694
rect 224622 657458 224804 657694
rect 224204 621694 224804 657458
rect 224204 621458 224386 621694
rect 224622 621458 224804 621694
rect 224204 585694 224804 621458
rect 224204 585458 224386 585694
rect 224622 585458 224804 585694
rect 224204 549694 224804 585458
rect 224204 549458 224386 549694
rect 224622 549458 224804 549694
rect 224204 513694 224804 549458
rect 224204 513458 224386 513694
rect 224622 513458 224804 513694
rect 224204 477694 224804 513458
rect 224204 477458 224386 477694
rect 224622 477458 224804 477694
rect 224204 441694 224804 477458
rect 224204 441458 224386 441694
rect 224622 441458 224804 441694
rect 224204 405694 224804 441458
rect 224204 405458 224386 405694
rect 224622 405458 224804 405694
rect 224204 369694 224804 405458
rect 224204 369458 224386 369694
rect 224622 369458 224804 369694
rect 224204 333694 224804 369458
rect 224204 333458 224386 333694
rect 224622 333458 224804 333694
rect 224204 297694 224804 333458
rect 224204 297458 224386 297694
rect 224622 297458 224804 297694
rect 224204 261694 224804 297458
rect 224204 261458 224386 261694
rect 224622 261458 224804 261694
rect 224204 242304 224804 261458
rect 227904 697394 228504 710042
rect 245904 711558 246504 711590
rect 245904 711322 246086 711558
rect 246322 711322 246504 711558
rect 245904 711238 246504 711322
rect 245904 711002 246086 711238
rect 246322 711002 246504 711238
rect 242204 709638 242804 709670
rect 242204 709402 242386 709638
rect 242622 709402 242804 709638
rect 242204 709318 242804 709402
rect 242204 709082 242386 709318
rect 242622 709082 242804 709318
rect 238504 707718 239104 707750
rect 238504 707482 238686 707718
rect 238922 707482 239104 707718
rect 238504 707398 239104 707482
rect 238504 707162 238686 707398
rect 238922 707162 239104 707398
rect 227904 697158 228086 697394
rect 228322 697158 228504 697394
rect 227904 661394 228504 697158
rect 227904 661158 228086 661394
rect 228322 661158 228504 661394
rect 227904 625394 228504 661158
rect 227904 625158 228086 625394
rect 228322 625158 228504 625394
rect 227904 589394 228504 625158
rect 227904 589158 228086 589394
rect 228322 589158 228504 589394
rect 227904 553394 228504 589158
rect 227904 553158 228086 553394
rect 228322 553158 228504 553394
rect 227904 517394 228504 553158
rect 227904 517158 228086 517394
rect 228322 517158 228504 517394
rect 227904 481394 228504 517158
rect 227904 481158 228086 481394
rect 228322 481158 228504 481394
rect 227904 445394 228504 481158
rect 227904 445158 228086 445394
rect 228322 445158 228504 445394
rect 227904 409394 228504 445158
rect 227904 409158 228086 409394
rect 228322 409158 228504 409394
rect 227904 373394 228504 409158
rect 227904 373158 228086 373394
rect 228322 373158 228504 373394
rect 227904 337394 228504 373158
rect 234804 705798 235404 705830
rect 234804 705562 234986 705798
rect 235222 705562 235404 705798
rect 234804 705478 235404 705562
rect 234804 705242 234986 705478
rect 235222 705242 235404 705478
rect 234804 668294 235404 705242
rect 234804 668058 234986 668294
rect 235222 668058 235404 668294
rect 234804 632294 235404 668058
rect 234804 632058 234986 632294
rect 235222 632058 235404 632294
rect 234804 596294 235404 632058
rect 234804 596058 234986 596294
rect 235222 596058 235404 596294
rect 234804 560294 235404 596058
rect 234804 560058 234986 560294
rect 235222 560058 235404 560294
rect 234804 524294 235404 560058
rect 234804 524058 234986 524294
rect 235222 524058 235404 524294
rect 234804 488294 235404 524058
rect 234804 488058 234986 488294
rect 235222 488058 235404 488294
rect 234804 452294 235404 488058
rect 234804 452058 234986 452294
rect 235222 452058 235404 452294
rect 234804 416294 235404 452058
rect 234804 416058 234986 416294
rect 235222 416058 235404 416294
rect 234804 380294 235404 416058
rect 234804 380058 234986 380294
rect 235222 380058 235404 380294
rect 234804 344294 235404 380058
rect 234804 344058 234986 344294
rect 235222 344058 235404 344294
rect 233187 337652 233253 337653
rect 233187 337588 233188 337652
rect 233252 337588 233253 337652
rect 233187 337587 233253 337588
rect 231899 337516 231965 337517
rect 231899 337452 231900 337516
rect 231964 337452 231965 337516
rect 231899 337451 231965 337452
rect 227904 337158 228086 337394
rect 228322 337158 228504 337394
rect 227904 301394 228504 337158
rect 227904 301158 228086 301394
rect 228322 301158 228504 301394
rect 227904 265394 228504 301158
rect 227904 265158 228086 265394
rect 228322 265158 228504 265394
rect 227904 242304 228504 265158
rect 59123 239732 59189 239733
rect 59123 239668 59124 239732
rect 59188 239668 59189 239732
rect 59123 239667 59189 239668
rect 75867 239732 75933 239733
rect 75867 239668 75868 239732
rect 75932 239668 75933 239732
rect 75867 239667 75933 239668
rect 58203 39948 58269 39949
rect 58203 39884 58204 39948
rect 58268 39884 58269 39948
rect 58203 39883 58269 39884
rect 59126 38317 59186 239667
rect 59307 239460 59373 239461
rect 59307 239396 59308 239460
rect 59372 239396 59373 239460
rect 59307 239395 59373 239396
rect 59123 38316 59189 38317
rect 59123 38252 59124 38316
rect 59188 38252 59189 38316
rect 59123 38251 59189 38252
rect 59310 38181 59370 239395
rect 59568 236294 59888 236476
rect 59568 236058 59610 236294
rect 59846 236058 59888 236294
rect 59568 235876 59888 236058
rect 90288 236294 90608 236476
rect 90288 236058 90330 236294
rect 90566 236058 90608 236294
rect 90288 235876 90608 236058
rect 121008 236294 121328 236476
rect 121008 236058 121050 236294
rect 121286 236058 121328 236294
rect 121008 235876 121328 236058
rect 151728 236294 152048 236476
rect 151728 236058 151770 236294
rect 152006 236058 152048 236294
rect 151728 235876 152048 236058
rect 182448 236294 182768 236476
rect 182448 236058 182490 236294
rect 182726 236058 182768 236294
rect 182448 235876 182768 236058
rect 213168 236294 213488 236476
rect 213168 236058 213210 236294
rect 213446 236058 213488 236294
rect 213168 235876 213488 236058
rect 74928 218294 75248 218476
rect 74928 218058 74970 218294
rect 75206 218058 75248 218294
rect 74928 217876 75248 218058
rect 105648 218294 105968 218476
rect 105648 218058 105690 218294
rect 105926 218058 105968 218294
rect 105648 217876 105968 218058
rect 136368 218294 136688 218476
rect 136368 218058 136410 218294
rect 136646 218058 136688 218294
rect 136368 217876 136688 218058
rect 167088 218294 167408 218476
rect 167088 218058 167130 218294
rect 167366 218058 167408 218294
rect 167088 217876 167408 218058
rect 197808 218294 198128 218476
rect 197808 218058 197850 218294
rect 198086 218058 198128 218294
rect 197808 217876 198128 218058
rect 228528 218294 228848 218476
rect 228528 218058 228570 218294
rect 228806 218058 228848 218294
rect 228528 217876 228848 218058
rect 59568 200294 59888 200476
rect 59568 200058 59610 200294
rect 59846 200058 59888 200294
rect 59568 199876 59888 200058
rect 90288 200294 90608 200476
rect 90288 200058 90330 200294
rect 90566 200058 90608 200294
rect 90288 199876 90608 200058
rect 121008 200294 121328 200476
rect 121008 200058 121050 200294
rect 121286 200058 121328 200294
rect 121008 199876 121328 200058
rect 151728 200294 152048 200476
rect 151728 200058 151770 200294
rect 152006 200058 152048 200294
rect 151728 199876 152048 200058
rect 182448 200294 182768 200476
rect 182448 200058 182490 200294
rect 182726 200058 182768 200294
rect 182448 199876 182768 200058
rect 213168 200294 213488 200476
rect 213168 200058 213210 200294
rect 213446 200058 213488 200294
rect 213168 199876 213488 200058
rect 74928 182294 75248 182476
rect 74928 182058 74970 182294
rect 75206 182058 75248 182294
rect 74928 181876 75248 182058
rect 105648 182294 105968 182476
rect 105648 182058 105690 182294
rect 105926 182058 105968 182294
rect 105648 181876 105968 182058
rect 136368 182294 136688 182476
rect 136368 182058 136410 182294
rect 136646 182058 136688 182294
rect 136368 181876 136688 182058
rect 167088 182294 167408 182476
rect 167088 182058 167130 182294
rect 167366 182058 167408 182294
rect 167088 181876 167408 182058
rect 197808 182294 198128 182476
rect 197808 182058 197850 182294
rect 198086 182058 198128 182294
rect 197808 181876 198128 182058
rect 228528 182294 228848 182476
rect 228528 182058 228570 182294
rect 228806 182058 228848 182294
rect 228528 181876 228848 182058
rect 59568 164294 59888 164476
rect 59568 164058 59610 164294
rect 59846 164058 59888 164294
rect 59568 163876 59888 164058
rect 90288 164294 90608 164476
rect 90288 164058 90330 164294
rect 90566 164058 90608 164294
rect 90288 163876 90608 164058
rect 121008 164294 121328 164476
rect 121008 164058 121050 164294
rect 121286 164058 121328 164294
rect 121008 163876 121328 164058
rect 151728 164294 152048 164476
rect 151728 164058 151770 164294
rect 152006 164058 152048 164294
rect 151728 163876 152048 164058
rect 182448 164294 182768 164476
rect 182448 164058 182490 164294
rect 182726 164058 182768 164294
rect 182448 163876 182768 164058
rect 213168 164294 213488 164476
rect 213168 164058 213210 164294
rect 213446 164058 213488 164294
rect 213168 163876 213488 164058
rect 74928 146294 75248 146476
rect 74928 146058 74970 146294
rect 75206 146058 75248 146294
rect 74928 145876 75248 146058
rect 105648 146294 105968 146476
rect 105648 146058 105690 146294
rect 105926 146058 105968 146294
rect 105648 145876 105968 146058
rect 136368 146294 136688 146476
rect 136368 146058 136410 146294
rect 136646 146058 136688 146294
rect 136368 145876 136688 146058
rect 167088 146294 167408 146476
rect 167088 146058 167130 146294
rect 167366 146058 167408 146294
rect 167088 145876 167408 146058
rect 197808 146294 198128 146476
rect 197808 146058 197850 146294
rect 198086 146058 198128 146294
rect 197808 145876 198128 146058
rect 228528 146294 228848 146476
rect 228528 146058 228570 146294
rect 228806 146058 228848 146294
rect 228528 145876 228848 146058
rect 59568 128294 59888 128476
rect 59568 128058 59610 128294
rect 59846 128058 59888 128294
rect 59568 127876 59888 128058
rect 90288 128294 90608 128476
rect 90288 128058 90330 128294
rect 90566 128058 90608 128294
rect 90288 127876 90608 128058
rect 121008 128294 121328 128476
rect 121008 128058 121050 128294
rect 121286 128058 121328 128294
rect 121008 127876 121328 128058
rect 151728 128294 152048 128476
rect 151728 128058 151770 128294
rect 152006 128058 152048 128294
rect 151728 127876 152048 128058
rect 182448 128294 182768 128476
rect 182448 128058 182490 128294
rect 182726 128058 182768 128294
rect 182448 127876 182768 128058
rect 213168 128294 213488 128476
rect 213168 128058 213210 128294
rect 213446 128058 213488 128294
rect 213168 127876 213488 128058
rect 74928 110294 75248 110476
rect 74928 110058 74970 110294
rect 75206 110058 75248 110294
rect 74928 109876 75248 110058
rect 105648 110294 105968 110476
rect 105648 110058 105690 110294
rect 105926 110058 105968 110294
rect 105648 109876 105968 110058
rect 136368 110294 136688 110476
rect 136368 110058 136410 110294
rect 136646 110058 136688 110294
rect 136368 109876 136688 110058
rect 167088 110294 167408 110476
rect 167088 110058 167130 110294
rect 167366 110058 167408 110294
rect 167088 109876 167408 110058
rect 197808 110294 198128 110476
rect 197808 110058 197850 110294
rect 198086 110058 198128 110294
rect 197808 109876 198128 110058
rect 228528 110294 228848 110476
rect 228528 110058 228570 110294
rect 228806 110058 228848 110294
rect 228528 109876 228848 110058
rect 59568 92294 59888 92476
rect 59568 92058 59610 92294
rect 59846 92058 59888 92294
rect 59568 91876 59888 92058
rect 90288 92294 90608 92476
rect 90288 92058 90330 92294
rect 90566 92058 90608 92294
rect 90288 91876 90608 92058
rect 121008 92294 121328 92476
rect 121008 92058 121050 92294
rect 121286 92058 121328 92294
rect 121008 91876 121328 92058
rect 151728 92294 152048 92476
rect 151728 92058 151770 92294
rect 152006 92058 152048 92294
rect 151728 91876 152048 92058
rect 182448 92294 182768 92476
rect 182448 92058 182490 92294
rect 182726 92058 182768 92294
rect 182448 91876 182768 92058
rect 213168 92294 213488 92476
rect 213168 92058 213210 92294
rect 213446 92058 213488 92294
rect 213168 91876 213488 92058
rect 74928 74294 75248 74476
rect 74928 74058 74970 74294
rect 75206 74058 75248 74294
rect 74928 73876 75248 74058
rect 105648 74294 105968 74476
rect 105648 74058 105690 74294
rect 105926 74058 105968 74294
rect 105648 73876 105968 74058
rect 136368 74294 136688 74476
rect 136368 74058 136410 74294
rect 136646 74058 136688 74294
rect 136368 73876 136688 74058
rect 167088 74294 167408 74476
rect 167088 74058 167130 74294
rect 167366 74058 167408 74294
rect 167088 73876 167408 74058
rect 197808 74294 198128 74476
rect 197808 74058 197850 74294
rect 198086 74058 198128 74294
rect 197808 73876 198128 74058
rect 228528 74294 228848 74476
rect 228528 74058 228570 74294
rect 228806 74058 228848 74294
rect 228528 73876 228848 74058
rect 59568 56294 59888 56476
rect 59568 56058 59610 56294
rect 59846 56058 59888 56294
rect 59568 55876 59888 56058
rect 90288 56294 90608 56476
rect 90288 56058 90330 56294
rect 90566 56058 90608 56294
rect 90288 55876 90608 56058
rect 121008 56294 121328 56476
rect 121008 56058 121050 56294
rect 121286 56058 121328 56294
rect 121008 55876 121328 56058
rect 151728 56294 152048 56476
rect 151728 56058 151770 56294
rect 152006 56058 152048 56294
rect 151728 55876 152048 56058
rect 182448 56294 182768 56476
rect 182448 56058 182490 56294
rect 182726 56058 182768 56294
rect 182448 55876 182768 56058
rect 213168 56294 213488 56476
rect 213168 56058 213210 56294
rect 213446 56058 213488 56294
rect 213168 55876 213488 56058
rect 231902 38453 231962 337451
rect 233190 38589 233250 337587
rect 234804 308294 235404 344058
rect 234804 308058 234986 308294
rect 235222 308058 235404 308294
rect 234804 272294 235404 308058
rect 234804 272058 234986 272294
rect 235222 272058 235404 272294
rect 234804 242304 235404 272058
rect 238504 671994 239104 707162
rect 238504 671758 238686 671994
rect 238922 671758 239104 671994
rect 238504 635994 239104 671758
rect 238504 635758 238686 635994
rect 238922 635758 239104 635994
rect 238504 599994 239104 635758
rect 238504 599758 238686 599994
rect 238922 599758 239104 599994
rect 238504 563994 239104 599758
rect 238504 563758 238686 563994
rect 238922 563758 239104 563994
rect 238504 527994 239104 563758
rect 238504 527758 238686 527994
rect 238922 527758 239104 527994
rect 238504 491994 239104 527758
rect 238504 491758 238686 491994
rect 238922 491758 239104 491994
rect 238504 455994 239104 491758
rect 238504 455758 238686 455994
rect 238922 455758 239104 455994
rect 238504 419994 239104 455758
rect 238504 419758 238686 419994
rect 238922 419758 239104 419994
rect 238504 383994 239104 419758
rect 238504 383758 238686 383994
rect 238922 383758 239104 383994
rect 238504 347994 239104 383758
rect 238504 347758 238686 347994
rect 238922 347758 239104 347994
rect 238504 311994 239104 347758
rect 238504 311758 238686 311994
rect 238922 311758 239104 311994
rect 238504 275994 239104 311758
rect 238504 275758 238686 275994
rect 238922 275758 239104 275994
rect 238504 242304 239104 275758
rect 242204 675694 242804 709082
rect 242204 675458 242386 675694
rect 242622 675458 242804 675694
rect 242204 639694 242804 675458
rect 242204 639458 242386 639694
rect 242622 639458 242804 639694
rect 242204 603694 242804 639458
rect 242204 603458 242386 603694
rect 242622 603458 242804 603694
rect 242204 567694 242804 603458
rect 242204 567458 242386 567694
rect 242622 567458 242804 567694
rect 242204 531694 242804 567458
rect 242204 531458 242386 531694
rect 242622 531458 242804 531694
rect 242204 495694 242804 531458
rect 242204 495458 242386 495694
rect 242622 495458 242804 495694
rect 242204 459694 242804 495458
rect 242204 459458 242386 459694
rect 242622 459458 242804 459694
rect 242204 423694 242804 459458
rect 242204 423458 242386 423694
rect 242622 423458 242804 423694
rect 242204 387694 242804 423458
rect 242204 387458 242386 387694
rect 242622 387458 242804 387694
rect 242204 351694 242804 387458
rect 242204 351458 242386 351694
rect 242622 351458 242804 351694
rect 242204 315694 242804 351458
rect 242204 315458 242386 315694
rect 242622 315458 242804 315694
rect 242204 279694 242804 315458
rect 242204 279458 242386 279694
rect 242622 279458 242804 279694
rect 242204 243694 242804 279458
rect 242204 243458 242386 243694
rect 242622 243458 242804 243694
rect 242204 207694 242804 243458
rect 242204 207458 242386 207694
rect 242622 207458 242804 207694
rect 242204 171694 242804 207458
rect 242204 171458 242386 171694
rect 242622 171458 242804 171694
rect 242204 135694 242804 171458
rect 242204 135458 242386 135694
rect 242622 135458 242804 135694
rect 242204 99694 242804 135458
rect 242204 99458 242386 99694
rect 242622 99458 242804 99694
rect 242204 63694 242804 99458
rect 242204 63458 242386 63694
rect 242622 63458 242804 63694
rect 233187 38588 233253 38589
rect 233187 38524 233188 38588
rect 233252 38524 233253 38588
rect 233187 38523 233253 38524
rect 231899 38452 231965 38453
rect 231899 38388 231900 38452
rect 231964 38388 231965 38452
rect 231899 38387 231965 38388
rect 59307 38180 59373 38181
rect 59307 38116 59308 38180
rect 59372 38116 59373 38180
rect 59307 38115 59373 38116
rect 57835 37772 57901 37773
rect 57835 37708 57836 37772
rect 57900 37708 57901 37772
rect 57835 37707 57901 37708
rect 54804 20058 54986 20294
rect 55222 20058 55404 20294
rect 54804 -1306 55404 20058
rect 54804 -1542 54986 -1306
rect 55222 -1542 55404 -1306
rect 54804 -1626 55404 -1542
rect 54804 -1862 54986 -1626
rect 55222 -1862 55404 -1626
rect 54804 -1894 55404 -1862
rect 58504 23994 59104 38000
rect 58504 23758 58686 23994
rect 58922 23758 59104 23994
rect 58504 -3226 59104 23758
rect 58504 -3462 58686 -3226
rect 58922 -3462 59104 -3226
rect 58504 -3546 59104 -3462
rect 58504 -3782 58686 -3546
rect 58922 -3782 59104 -3546
rect 58504 -3814 59104 -3782
rect 62204 27694 62804 38000
rect 62204 27458 62386 27694
rect 62622 27458 62804 27694
rect 62204 -5146 62804 27458
rect 62204 -5382 62386 -5146
rect 62622 -5382 62804 -5146
rect 62204 -5466 62804 -5382
rect 62204 -5702 62386 -5466
rect 62622 -5702 62804 -5466
rect 62204 -5734 62804 -5702
rect 65904 31394 66504 38000
rect 65904 31158 66086 31394
rect 66322 31158 66504 31394
rect 47904 -6342 48086 -6106
rect 48322 -6342 48504 -6106
rect 47904 -6426 48504 -6342
rect 47904 -6662 48086 -6426
rect 48322 -6662 48504 -6426
rect 47904 -7654 48504 -6662
rect 65904 -7066 66504 31158
rect 72804 2294 73404 38000
rect 72804 2058 72986 2294
rect 73222 2058 73404 2294
rect 72804 -346 73404 2058
rect 72804 -582 72986 -346
rect 73222 -582 73404 -346
rect 72804 -666 73404 -582
rect 72804 -902 72986 -666
rect 73222 -902 73404 -666
rect 72804 -1894 73404 -902
rect 76504 5994 77104 38000
rect 76504 5758 76686 5994
rect 76922 5758 77104 5994
rect 76504 -2266 77104 5758
rect 76504 -2502 76686 -2266
rect 76922 -2502 77104 -2266
rect 76504 -2586 77104 -2502
rect 76504 -2822 76686 -2586
rect 76922 -2822 77104 -2586
rect 76504 -3814 77104 -2822
rect 80204 9694 80804 38000
rect 80204 9458 80386 9694
rect 80622 9458 80804 9694
rect 80204 -4186 80804 9458
rect 80204 -4422 80386 -4186
rect 80622 -4422 80804 -4186
rect 80204 -4506 80804 -4422
rect 80204 -4742 80386 -4506
rect 80622 -4742 80804 -4506
rect 80204 -5734 80804 -4742
rect 83904 13394 84504 38000
rect 83904 13158 84086 13394
rect 84322 13158 84504 13394
rect 65904 -7302 66086 -7066
rect 66322 -7302 66504 -7066
rect 65904 -7386 66504 -7302
rect 65904 -7622 66086 -7386
rect 66322 -7622 66504 -7386
rect 65904 -7654 66504 -7622
rect 83904 -6106 84504 13158
rect 90804 20294 91404 38000
rect 90804 20058 90986 20294
rect 91222 20058 91404 20294
rect 90804 -1306 91404 20058
rect 90804 -1542 90986 -1306
rect 91222 -1542 91404 -1306
rect 90804 -1626 91404 -1542
rect 90804 -1862 90986 -1626
rect 91222 -1862 91404 -1626
rect 90804 -1894 91404 -1862
rect 94504 23994 95104 38000
rect 94504 23758 94686 23994
rect 94922 23758 95104 23994
rect 94504 -3226 95104 23758
rect 94504 -3462 94686 -3226
rect 94922 -3462 95104 -3226
rect 94504 -3546 95104 -3462
rect 94504 -3782 94686 -3546
rect 94922 -3782 95104 -3546
rect 94504 -3814 95104 -3782
rect 98204 27694 98804 38000
rect 98204 27458 98386 27694
rect 98622 27458 98804 27694
rect 98204 -5146 98804 27458
rect 98204 -5382 98386 -5146
rect 98622 -5382 98804 -5146
rect 98204 -5466 98804 -5382
rect 98204 -5702 98386 -5466
rect 98622 -5702 98804 -5466
rect 98204 -5734 98804 -5702
rect 101904 31394 102504 38000
rect 101904 31158 102086 31394
rect 102322 31158 102504 31394
rect 83904 -6342 84086 -6106
rect 84322 -6342 84504 -6106
rect 83904 -6426 84504 -6342
rect 83904 -6662 84086 -6426
rect 84322 -6662 84504 -6426
rect 83904 -7654 84504 -6662
rect 101904 -7066 102504 31158
rect 108804 2294 109404 38000
rect 108804 2058 108986 2294
rect 109222 2058 109404 2294
rect 108804 -346 109404 2058
rect 108804 -582 108986 -346
rect 109222 -582 109404 -346
rect 108804 -666 109404 -582
rect 108804 -902 108986 -666
rect 109222 -902 109404 -666
rect 108804 -1894 109404 -902
rect 112504 5994 113104 38000
rect 112504 5758 112686 5994
rect 112922 5758 113104 5994
rect 112504 -2266 113104 5758
rect 112504 -2502 112686 -2266
rect 112922 -2502 113104 -2266
rect 112504 -2586 113104 -2502
rect 112504 -2822 112686 -2586
rect 112922 -2822 113104 -2586
rect 112504 -3814 113104 -2822
rect 116204 9694 116804 38000
rect 116204 9458 116386 9694
rect 116622 9458 116804 9694
rect 116204 -4186 116804 9458
rect 116204 -4422 116386 -4186
rect 116622 -4422 116804 -4186
rect 116204 -4506 116804 -4422
rect 116204 -4742 116386 -4506
rect 116622 -4742 116804 -4506
rect 116204 -5734 116804 -4742
rect 119904 13394 120504 38000
rect 119904 13158 120086 13394
rect 120322 13158 120504 13394
rect 101904 -7302 102086 -7066
rect 102322 -7302 102504 -7066
rect 101904 -7386 102504 -7302
rect 101904 -7622 102086 -7386
rect 102322 -7622 102504 -7386
rect 101904 -7654 102504 -7622
rect 119904 -6106 120504 13158
rect 126804 20294 127404 38000
rect 126804 20058 126986 20294
rect 127222 20058 127404 20294
rect 126804 -1306 127404 20058
rect 126804 -1542 126986 -1306
rect 127222 -1542 127404 -1306
rect 126804 -1626 127404 -1542
rect 126804 -1862 126986 -1626
rect 127222 -1862 127404 -1626
rect 126804 -1894 127404 -1862
rect 130504 23994 131104 38000
rect 130504 23758 130686 23994
rect 130922 23758 131104 23994
rect 130504 -3226 131104 23758
rect 130504 -3462 130686 -3226
rect 130922 -3462 131104 -3226
rect 130504 -3546 131104 -3462
rect 130504 -3782 130686 -3546
rect 130922 -3782 131104 -3546
rect 130504 -3814 131104 -3782
rect 134204 27694 134804 38000
rect 134204 27458 134386 27694
rect 134622 27458 134804 27694
rect 134204 -5146 134804 27458
rect 134204 -5382 134386 -5146
rect 134622 -5382 134804 -5146
rect 134204 -5466 134804 -5382
rect 134204 -5702 134386 -5466
rect 134622 -5702 134804 -5466
rect 134204 -5734 134804 -5702
rect 137904 31394 138504 38000
rect 137904 31158 138086 31394
rect 138322 31158 138504 31394
rect 119904 -6342 120086 -6106
rect 120322 -6342 120504 -6106
rect 119904 -6426 120504 -6342
rect 119904 -6662 120086 -6426
rect 120322 -6662 120504 -6426
rect 119904 -7654 120504 -6662
rect 137904 -7066 138504 31158
rect 144804 2294 145404 38000
rect 144804 2058 144986 2294
rect 145222 2058 145404 2294
rect 144804 -346 145404 2058
rect 144804 -582 144986 -346
rect 145222 -582 145404 -346
rect 144804 -666 145404 -582
rect 144804 -902 144986 -666
rect 145222 -902 145404 -666
rect 144804 -1894 145404 -902
rect 148504 5994 149104 38000
rect 148504 5758 148686 5994
rect 148922 5758 149104 5994
rect 148504 -2266 149104 5758
rect 148504 -2502 148686 -2266
rect 148922 -2502 149104 -2266
rect 148504 -2586 149104 -2502
rect 148504 -2822 148686 -2586
rect 148922 -2822 149104 -2586
rect 148504 -3814 149104 -2822
rect 152204 9694 152804 38000
rect 152204 9458 152386 9694
rect 152622 9458 152804 9694
rect 152204 -4186 152804 9458
rect 152204 -4422 152386 -4186
rect 152622 -4422 152804 -4186
rect 152204 -4506 152804 -4422
rect 152204 -4742 152386 -4506
rect 152622 -4742 152804 -4506
rect 152204 -5734 152804 -4742
rect 155904 13394 156504 38000
rect 155904 13158 156086 13394
rect 156322 13158 156504 13394
rect 137904 -7302 138086 -7066
rect 138322 -7302 138504 -7066
rect 137904 -7386 138504 -7302
rect 137904 -7622 138086 -7386
rect 138322 -7622 138504 -7386
rect 137904 -7654 138504 -7622
rect 155904 -6106 156504 13158
rect 162804 20294 163404 38000
rect 162804 20058 162986 20294
rect 163222 20058 163404 20294
rect 162804 -1306 163404 20058
rect 162804 -1542 162986 -1306
rect 163222 -1542 163404 -1306
rect 162804 -1626 163404 -1542
rect 162804 -1862 162986 -1626
rect 163222 -1862 163404 -1626
rect 162804 -1894 163404 -1862
rect 166504 23994 167104 38000
rect 166504 23758 166686 23994
rect 166922 23758 167104 23994
rect 166504 -3226 167104 23758
rect 166504 -3462 166686 -3226
rect 166922 -3462 167104 -3226
rect 166504 -3546 167104 -3462
rect 166504 -3782 166686 -3546
rect 166922 -3782 167104 -3546
rect 166504 -3814 167104 -3782
rect 170204 27694 170804 38000
rect 170204 27458 170386 27694
rect 170622 27458 170804 27694
rect 170204 -5146 170804 27458
rect 170204 -5382 170386 -5146
rect 170622 -5382 170804 -5146
rect 170204 -5466 170804 -5382
rect 170204 -5702 170386 -5466
rect 170622 -5702 170804 -5466
rect 170204 -5734 170804 -5702
rect 173904 31394 174504 38000
rect 173904 31158 174086 31394
rect 174322 31158 174504 31394
rect 155904 -6342 156086 -6106
rect 156322 -6342 156504 -6106
rect 155904 -6426 156504 -6342
rect 155904 -6662 156086 -6426
rect 156322 -6662 156504 -6426
rect 155904 -7654 156504 -6662
rect 173904 -7066 174504 31158
rect 180804 2294 181404 38000
rect 180804 2058 180986 2294
rect 181222 2058 181404 2294
rect 180804 -346 181404 2058
rect 180804 -582 180986 -346
rect 181222 -582 181404 -346
rect 180804 -666 181404 -582
rect 180804 -902 180986 -666
rect 181222 -902 181404 -666
rect 180804 -1894 181404 -902
rect 184504 5994 185104 38000
rect 184504 5758 184686 5994
rect 184922 5758 185104 5994
rect 184504 -2266 185104 5758
rect 184504 -2502 184686 -2266
rect 184922 -2502 185104 -2266
rect 184504 -2586 185104 -2502
rect 184504 -2822 184686 -2586
rect 184922 -2822 185104 -2586
rect 184504 -3814 185104 -2822
rect 188204 9694 188804 38000
rect 188204 9458 188386 9694
rect 188622 9458 188804 9694
rect 188204 -4186 188804 9458
rect 188204 -4422 188386 -4186
rect 188622 -4422 188804 -4186
rect 188204 -4506 188804 -4422
rect 188204 -4742 188386 -4506
rect 188622 -4742 188804 -4506
rect 188204 -5734 188804 -4742
rect 191904 13394 192504 38000
rect 191904 13158 192086 13394
rect 192322 13158 192504 13394
rect 173904 -7302 174086 -7066
rect 174322 -7302 174504 -7066
rect 173904 -7386 174504 -7302
rect 173904 -7622 174086 -7386
rect 174322 -7622 174504 -7386
rect 173904 -7654 174504 -7622
rect 191904 -6106 192504 13158
rect 198804 20294 199404 38000
rect 198804 20058 198986 20294
rect 199222 20058 199404 20294
rect 198804 -1306 199404 20058
rect 198804 -1542 198986 -1306
rect 199222 -1542 199404 -1306
rect 198804 -1626 199404 -1542
rect 198804 -1862 198986 -1626
rect 199222 -1862 199404 -1626
rect 198804 -1894 199404 -1862
rect 202504 23994 203104 38000
rect 202504 23758 202686 23994
rect 202922 23758 203104 23994
rect 202504 -3226 203104 23758
rect 202504 -3462 202686 -3226
rect 202922 -3462 203104 -3226
rect 202504 -3546 203104 -3462
rect 202504 -3782 202686 -3546
rect 202922 -3782 203104 -3546
rect 202504 -3814 203104 -3782
rect 206204 27694 206804 38000
rect 206204 27458 206386 27694
rect 206622 27458 206804 27694
rect 206204 -5146 206804 27458
rect 206204 -5382 206386 -5146
rect 206622 -5382 206804 -5146
rect 206204 -5466 206804 -5382
rect 206204 -5702 206386 -5466
rect 206622 -5702 206804 -5466
rect 206204 -5734 206804 -5702
rect 209904 31394 210504 38000
rect 209904 31158 210086 31394
rect 210322 31158 210504 31394
rect 191904 -6342 192086 -6106
rect 192322 -6342 192504 -6106
rect 191904 -6426 192504 -6342
rect 191904 -6662 192086 -6426
rect 192322 -6662 192504 -6426
rect 191904 -7654 192504 -6662
rect 209904 -7066 210504 31158
rect 216804 2294 217404 38000
rect 216804 2058 216986 2294
rect 217222 2058 217404 2294
rect 216804 -346 217404 2058
rect 216804 -582 216986 -346
rect 217222 -582 217404 -346
rect 216804 -666 217404 -582
rect 216804 -902 216986 -666
rect 217222 -902 217404 -666
rect 216804 -1894 217404 -902
rect 220504 5994 221104 38000
rect 220504 5758 220686 5994
rect 220922 5758 221104 5994
rect 220504 -2266 221104 5758
rect 220504 -2502 220686 -2266
rect 220922 -2502 221104 -2266
rect 220504 -2586 221104 -2502
rect 220504 -2822 220686 -2586
rect 220922 -2822 221104 -2586
rect 220504 -3814 221104 -2822
rect 224204 9694 224804 38000
rect 224204 9458 224386 9694
rect 224622 9458 224804 9694
rect 224204 -4186 224804 9458
rect 224204 -4422 224386 -4186
rect 224622 -4422 224804 -4186
rect 224204 -4506 224804 -4422
rect 224204 -4742 224386 -4506
rect 224622 -4742 224804 -4506
rect 224204 -5734 224804 -4742
rect 227904 13394 228504 38000
rect 227904 13158 228086 13394
rect 228322 13158 228504 13394
rect 209904 -7302 210086 -7066
rect 210322 -7302 210504 -7066
rect 209904 -7386 210504 -7302
rect 209904 -7622 210086 -7386
rect 210322 -7622 210504 -7386
rect 209904 -7654 210504 -7622
rect 227904 -6106 228504 13158
rect 234804 20294 235404 38000
rect 234804 20058 234986 20294
rect 235222 20058 235404 20294
rect 234804 -1306 235404 20058
rect 234804 -1542 234986 -1306
rect 235222 -1542 235404 -1306
rect 234804 -1626 235404 -1542
rect 234804 -1862 234986 -1626
rect 235222 -1862 235404 -1626
rect 234804 -1894 235404 -1862
rect 238504 23994 239104 38000
rect 238504 23758 238686 23994
rect 238922 23758 239104 23994
rect 238504 -3226 239104 23758
rect 238504 -3462 238686 -3226
rect 238922 -3462 239104 -3226
rect 238504 -3546 239104 -3462
rect 238504 -3782 238686 -3546
rect 238922 -3782 239104 -3546
rect 238504 -3814 239104 -3782
rect 242204 27694 242804 63458
rect 242204 27458 242386 27694
rect 242622 27458 242804 27694
rect 242204 -5146 242804 27458
rect 242204 -5382 242386 -5146
rect 242622 -5382 242804 -5146
rect 242204 -5466 242804 -5382
rect 242204 -5702 242386 -5466
rect 242622 -5702 242804 -5466
rect 242204 -5734 242804 -5702
rect 245904 679394 246504 711002
rect 263904 710598 264504 711590
rect 263904 710362 264086 710598
rect 264322 710362 264504 710598
rect 263904 710278 264504 710362
rect 263904 710042 264086 710278
rect 264322 710042 264504 710278
rect 260204 708678 260804 709670
rect 260204 708442 260386 708678
rect 260622 708442 260804 708678
rect 260204 708358 260804 708442
rect 260204 708122 260386 708358
rect 260622 708122 260804 708358
rect 256504 706758 257104 707750
rect 256504 706522 256686 706758
rect 256922 706522 257104 706758
rect 256504 706438 257104 706522
rect 256504 706202 256686 706438
rect 256922 706202 257104 706438
rect 245904 679158 246086 679394
rect 246322 679158 246504 679394
rect 245904 643394 246504 679158
rect 245904 643158 246086 643394
rect 246322 643158 246504 643394
rect 245904 607394 246504 643158
rect 245904 607158 246086 607394
rect 246322 607158 246504 607394
rect 245904 571394 246504 607158
rect 245904 571158 246086 571394
rect 246322 571158 246504 571394
rect 245904 535394 246504 571158
rect 245904 535158 246086 535394
rect 246322 535158 246504 535394
rect 245904 499394 246504 535158
rect 245904 499158 246086 499394
rect 246322 499158 246504 499394
rect 245904 463394 246504 499158
rect 245904 463158 246086 463394
rect 246322 463158 246504 463394
rect 245904 427394 246504 463158
rect 245904 427158 246086 427394
rect 246322 427158 246504 427394
rect 245904 391394 246504 427158
rect 245904 391158 246086 391394
rect 246322 391158 246504 391394
rect 245904 355394 246504 391158
rect 245904 355158 246086 355394
rect 246322 355158 246504 355394
rect 245904 319394 246504 355158
rect 245904 319158 246086 319394
rect 246322 319158 246504 319394
rect 245904 283394 246504 319158
rect 245904 283158 246086 283394
rect 246322 283158 246504 283394
rect 245904 247394 246504 283158
rect 245904 247158 246086 247394
rect 246322 247158 246504 247394
rect 245904 211394 246504 247158
rect 245904 211158 246086 211394
rect 246322 211158 246504 211394
rect 245904 175394 246504 211158
rect 245904 175158 246086 175394
rect 246322 175158 246504 175394
rect 245904 139394 246504 175158
rect 245904 139158 246086 139394
rect 246322 139158 246504 139394
rect 245904 103394 246504 139158
rect 245904 103158 246086 103394
rect 246322 103158 246504 103394
rect 245904 67394 246504 103158
rect 245904 67158 246086 67394
rect 246322 67158 246504 67394
rect 245904 31394 246504 67158
rect 245904 31158 246086 31394
rect 246322 31158 246504 31394
rect 227904 -6342 228086 -6106
rect 228322 -6342 228504 -6106
rect 227904 -6426 228504 -6342
rect 227904 -6662 228086 -6426
rect 228322 -6662 228504 -6426
rect 227904 -7654 228504 -6662
rect 245904 -7066 246504 31158
rect 252804 704838 253404 705830
rect 252804 704602 252986 704838
rect 253222 704602 253404 704838
rect 252804 704518 253404 704602
rect 252804 704282 252986 704518
rect 253222 704282 253404 704518
rect 252804 686294 253404 704282
rect 252804 686058 252986 686294
rect 253222 686058 253404 686294
rect 252804 650294 253404 686058
rect 252804 650058 252986 650294
rect 253222 650058 253404 650294
rect 252804 614294 253404 650058
rect 252804 614058 252986 614294
rect 253222 614058 253404 614294
rect 252804 578294 253404 614058
rect 252804 578058 252986 578294
rect 253222 578058 253404 578294
rect 252804 542294 253404 578058
rect 252804 542058 252986 542294
rect 253222 542058 253404 542294
rect 252804 506294 253404 542058
rect 252804 506058 252986 506294
rect 253222 506058 253404 506294
rect 252804 470294 253404 506058
rect 252804 470058 252986 470294
rect 253222 470058 253404 470294
rect 252804 434294 253404 470058
rect 252804 434058 252986 434294
rect 253222 434058 253404 434294
rect 252804 398294 253404 434058
rect 252804 398058 252986 398294
rect 253222 398058 253404 398294
rect 252804 362294 253404 398058
rect 252804 362058 252986 362294
rect 253222 362058 253404 362294
rect 252804 326294 253404 362058
rect 252804 326058 252986 326294
rect 253222 326058 253404 326294
rect 252804 290294 253404 326058
rect 252804 290058 252986 290294
rect 253222 290058 253404 290294
rect 252804 254294 253404 290058
rect 252804 254058 252986 254294
rect 253222 254058 253404 254294
rect 252804 218294 253404 254058
rect 252804 218058 252986 218294
rect 253222 218058 253404 218294
rect 252804 182294 253404 218058
rect 252804 182058 252986 182294
rect 253222 182058 253404 182294
rect 252804 146294 253404 182058
rect 252804 146058 252986 146294
rect 253222 146058 253404 146294
rect 252804 110294 253404 146058
rect 252804 110058 252986 110294
rect 253222 110058 253404 110294
rect 252804 74294 253404 110058
rect 252804 74058 252986 74294
rect 253222 74058 253404 74294
rect 252804 38294 253404 74058
rect 252804 38058 252986 38294
rect 253222 38058 253404 38294
rect 252804 2294 253404 38058
rect 252804 2058 252986 2294
rect 253222 2058 253404 2294
rect 252804 -346 253404 2058
rect 252804 -582 252986 -346
rect 253222 -582 253404 -346
rect 252804 -666 253404 -582
rect 252804 -902 252986 -666
rect 253222 -902 253404 -666
rect 252804 -1894 253404 -902
rect 256504 689994 257104 706202
rect 256504 689758 256686 689994
rect 256922 689758 257104 689994
rect 256504 653994 257104 689758
rect 256504 653758 256686 653994
rect 256922 653758 257104 653994
rect 256504 617994 257104 653758
rect 256504 617758 256686 617994
rect 256922 617758 257104 617994
rect 256504 581994 257104 617758
rect 256504 581758 256686 581994
rect 256922 581758 257104 581994
rect 256504 545994 257104 581758
rect 256504 545758 256686 545994
rect 256922 545758 257104 545994
rect 256504 509994 257104 545758
rect 256504 509758 256686 509994
rect 256922 509758 257104 509994
rect 256504 473994 257104 509758
rect 256504 473758 256686 473994
rect 256922 473758 257104 473994
rect 256504 437994 257104 473758
rect 256504 437758 256686 437994
rect 256922 437758 257104 437994
rect 256504 401994 257104 437758
rect 256504 401758 256686 401994
rect 256922 401758 257104 401994
rect 256504 365994 257104 401758
rect 256504 365758 256686 365994
rect 256922 365758 257104 365994
rect 256504 329994 257104 365758
rect 256504 329758 256686 329994
rect 256922 329758 257104 329994
rect 256504 293994 257104 329758
rect 256504 293758 256686 293994
rect 256922 293758 257104 293994
rect 256504 257994 257104 293758
rect 256504 257758 256686 257994
rect 256922 257758 257104 257994
rect 256504 221994 257104 257758
rect 256504 221758 256686 221994
rect 256922 221758 257104 221994
rect 256504 185994 257104 221758
rect 256504 185758 256686 185994
rect 256922 185758 257104 185994
rect 256504 149994 257104 185758
rect 256504 149758 256686 149994
rect 256922 149758 257104 149994
rect 256504 113994 257104 149758
rect 256504 113758 256686 113994
rect 256922 113758 257104 113994
rect 256504 77994 257104 113758
rect 256504 77758 256686 77994
rect 256922 77758 257104 77994
rect 256504 41994 257104 77758
rect 256504 41758 256686 41994
rect 256922 41758 257104 41994
rect 256504 5994 257104 41758
rect 256504 5758 256686 5994
rect 256922 5758 257104 5994
rect 256504 -2266 257104 5758
rect 256504 -2502 256686 -2266
rect 256922 -2502 257104 -2266
rect 256504 -2586 257104 -2502
rect 256504 -2822 256686 -2586
rect 256922 -2822 257104 -2586
rect 256504 -3814 257104 -2822
rect 260204 693694 260804 708122
rect 260204 693458 260386 693694
rect 260622 693458 260804 693694
rect 260204 657694 260804 693458
rect 260204 657458 260386 657694
rect 260622 657458 260804 657694
rect 260204 621694 260804 657458
rect 260204 621458 260386 621694
rect 260622 621458 260804 621694
rect 260204 585694 260804 621458
rect 260204 585458 260386 585694
rect 260622 585458 260804 585694
rect 260204 549694 260804 585458
rect 260204 549458 260386 549694
rect 260622 549458 260804 549694
rect 260204 513694 260804 549458
rect 260204 513458 260386 513694
rect 260622 513458 260804 513694
rect 260204 477694 260804 513458
rect 260204 477458 260386 477694
rect 260622 477458 260804 477694
rect 260204 441694 260804 477458
rect 260204 441458 260386 441694
rect 260622 441458 260804 441694
rect 260204 405694 260804 441458
rect 260204 405458 260386 405694
rect 260622 405458 260804 405694
rect 260204 369694 260804 405458
rect 260204 369458 260386 369694
rect 260622 369458 260804 369694
rect 260204 333694 260804 369458
rect 260204 333458 260386 333694
rect 260622 333458 260804 333694
rect 260204 297694 260804 333458
rect 260204 297458 260386 297694
rect 260622 297458 260804 297694
rect 260204 261694 260804 297458
rect 260204 261458 260386 261694
rect 260622 261458 260804 261694
rect 260204 225694 260804 261458
rect 260204 225458 260386 225694
rect 260622 225458 260804 225694
rect 260204 189694 260804 225458
rect 260204 189458 260386 189694
rect 260622 189458 260804 189694
rect 260204 153694 260804 189458
rect 260204 153458 260386 153694
rect 260622 153458 260804 153694
rect 260204 117694 260804 153458
rect 260204 117458 260386 117694
rect 260622 117458 260804 117694
rect 260204 81694 260804 117458
rect 260204 81458 260386 81694
rect 260622 81458 260804 81694
rect 260204 45694 260804 81458
rect 260204 45458 260386 45694
rect 260622 45458 260804 45694
rect 260204 9694 260804 45458
rect 260204 9458 260386 9694
rect 260622 9458 260804 9694
rect 260204 -4186 260804 9458
rect 260204 -4422 260386 -4186
rect 260622 -4422 260804 -4186
rect 260204 -4506 260804 -4422
rect 260204 -4742 260386 -4506
rect 260622 -4742 260804 -4506
rect 260204 -5734 260804 -4742
rect 263904 697394 264504 710042
rect 281904 711558 282504 711590
rect 281904 711322 282086 711558
rect 282322 711322 282504 711558
rect 281904 711238 282504 711322
rect 281904 711002 282086 711238
rect 282322 711002 282504 711238
rect 278204 709638 278804 709670
rect 278204 709402 278386 709638
rect 278622 709402 278804 709638
rect 278204 709318 278804 709402
rect 278204 709082 278386 709318
rect 278622 709082 278804 709318
rect 274504 707718 275104 707750
rect 274504 707482 274686 707718
rect 274922 707482 275104 707718
rect 274504 707398 275104 707482
rect 274504 707162 274686 707398
rect 274922 707162 275104 707398
rect 263904 697158 264086 697394
rect 264322 697158 264504 697394
rect 263904 661394 264504 697158
rect 263904 661158 264086 661394
rect 264322 661158 264504 661394
rect 263904 625394 264504 661158
rect 263904 625158 264086 625394
rect 264322 625158 264504 625394
rect 263904 589394 264504 625158
rect 263904 589158 264086 589394
rect 264322 589158 264504 589394
rect 263904 553394 264504 589158
rect 263904 553158 264086 553394
rect 264322 553158 264504 553394
rect 263904 517394 264504 553158
rect 263904 517158 264086 517394
rect 264322 517158 264504 517394
rect 263904 481394 264504 517158
rect 263904 481158 264086 481394
rect 264322 481158 264504 481394
rect 263904 445394 264504 481158
rect 263904 445158 264086 445394
rect 264322 445158 264504 445394
rect 263904 409394 264504 445158
rect 263904 409158 264086 409394
rect 264322 409158 264504 409394
rect 263904 373394 264504 409158
rect 263904 373158 264086 373394
rect 264322 373158 264504 373394
rect 263904 337394 264504 373158
rect 263904 337158 264086 337394
rect 264322 337158 264504 337394
rect 263904 301394 264504 337158
rect 263904 301158 264086 301394
rect 264322 301158 264504 301394
rect 263904 265394 264504 301158
rect 263904 265158 264086 265394
rect 264322 265158 264504 265394
rect 263904 229394 264504 265158
rect 263904 229158 264086 229394
rect 264322 229158 264504 229394
rect 263904 193394 264504 229158
rect 263904 193158 264086 193394
rect 264322 193158 264504 193394
rect 263904 157394 264504 193158
rect 263904 157158 264086 157394
rect 264322 157158 264504 157394
rect 263904 121394 264504 157158
rect 263904 121158 264086 121394
rect 264322 121158 264504 121394
rect 263904 85394 264504 121158
rect 263904 85158 264086 85394
rect 264322 85158 264504 85394
rect 263904 49394 264504 85158
rect 263904 49158 264086 49394
rect 264322 49158 264504 49394
rect 263904 13394 264504 49158
rect 263904 13158 264086 13394
rect 264322 13158 264504 13394
rect 245904 -7302 246086 -7066
rect 246322 -7302 246504 -7066
rect 245904 -7386 246504 -7302
rect 245904 -7622 246086 -7386
rect 246322 -7622 246504 -7386
rect 245904 -7654 246504 -7622
rect 263904 -6106 264504 13158
rect 270804 705798 271404 705830
rect 270804 705562 270986 705798
rect 271222 705562 271404 705798
rect 270804 705478 271404 705562
rect 270804 705242 270986 705478
rect 271222 705242 271404 705478
rect 270804 668294 271404 705242
rect 270804 668058 270986 668294
rect 271222 668058 271404 668294
rect 270804 632294 271404 668058
rect 270804 632058 270986 632294
rect 271222 632058 271404 632294
rect 270804 596294 271404 632058
rect 270804 596058 270986 596294
rect 271222 596058 271404 596294
rect 270804 560294 271404 596058
rect 270804 560058 270986 560294
rect 271222 560058 271404 560294
rect 270804 524294 271404 560058
rect 270804 524058 270986 524294
rect 271222 524058 271404 524294
rect 270804 488294 271404 524058
rect 270804 488058 270986 488294
rect 271222 488058 271404 488294
rect 270804 452294 271404 488058
rect 270804 452058 270986 452294
rect 271222 452058 271404 452294
rect 270804 416294 271404 452058
rect 270804 416058 270986 416294
rect 271222 416058 271404 416294
rect 270804 380294 271404 416058
rect 270804 380058 270986 380294
rect 271222 380058 271404 380294
rect 270804 344294 271404 380058
rect 270804 344058 270986 344294
rect 271222 344058 271404 344294
rect 270804 308294 271404 344058
rect 270804 308058 270986 308294
rect 271222 308058 271404 308294
rect 270804 272294 271404 308058
rect 270804 272058 270986 272294
rect 271222 272058 271404 272294
rect 270804 236294 271404 272058
rect 270804 236058 270986 236294
rect 271222 236058 271404 236294
rect 270804 200294 271404 236058
rect 270804 200058 270986 200294
rect 271222 200058 271404 200294
rect 270804 164294 271404 200058
rect 270804 164058 270986 164294
rect 271222 164058 271404 164294
rect 270804 128294 271404 164058
rect 270804 128058 270986 128294
rect 271222 128058 271404 128294
rect 270804 92294 271404 128058
rect 270804 92058 270986 92294
rect 271222 92058 271404 92294
rect 270804 56294 271404 92058
rect 270804 56058 270986 56294
rect 271222 56058 271404 56294
rect 270804 20294 271404 56058
rect 270804 20058 270986 20294
rect 271222 20058 271404 20294
rect 270804 -1306 271404 20058
rect 270804 -1542 270986 -1306
rect 271222 -1542 271404 -1306
rect 270804 -1626 271404 -1542
rect 270804 -1862 270986 -1626
rect 271222 -1862 271404 -1626
rect 270804 -1894 271404 -1862
rect 274504 671994 275104 707162
rect 274504 671758 274686 671994
rect 274922 671758 275104 671994
rect 274504 635994 275104 671758
rect 274504 635758 274686 635994
rect 274922 635758 275104 635994
rect 274504 599994 275104 635758
rect 274504 599758 274686 599994
rect 274922 599758 275104 599994
rect 274504 563994 275104 599758
rect 274504 563758 274686 563994
rect 274922 563758 275104 563994
rect 274504 527994 275104 563758
rect 274504 527758 274686 527994
rect 274922 527758 275104 527994
rect 274504 491994 275104 527758
rect 274504 491758 274686 491994
rect 274922 491758 275104 491994
rect 274504 455994 275104 491758
rect 274504 455758 274686 455994
rect 274922 455758 275104 455994
rect 274504 419994 275104 455758
rect 274504 419758 274686 419994
rect 274922 419758 275104 419994
rect 274504 383994 275104 419758
rect 274504 383758 274686 383994
rect 274922 383758 275104 383994
rect 274504 347994 275104 383758
rect 274504 347758 274686 347994
rect 274922 347758 275104 347994
rect 274504 311994 275104 347758
rect 274504 311758 274686 311994
rect 274922 311758 275104 311994
rect 274504 275994 275104 311758
rect 274504 275758 274686 275994
rect 274922 275758 275104 275994
rect 274504 239994 275104 275758
rect 274504 239758 274686 239994
rect 274922 239758 275104 239994
rect 274504 203994 275104 239758
rect 274504 203758 274686 203994
rect 274922 203758 275104 203994
rect 274504 167994 275104 203758
rect 274504 167758 274686 167994
rect 274922 167758 275104 167994
rect 274504 131994 275104 167758
rect 274504 131758 274686 131994
rect 274922 131758 275104 131994
rect 274504 95994 275104 131758
rect 274504 95758 274686 95994
rect 274922 95758 275104 95994
rect 274504 59994 275104 95758
rect 274504 59758 274686 59994
rect 274922 59758 275104 59994
rect 274504 23994 275104 59758
rect 274504 23758 274686 23994
rect 274922 23758 275104 23994
rect 274504 -3226 275104 23758
rect 274504 -3462 274686 -3226
rect 274922 -3462 275104 -3226
rect 274504 -3546 275104 -3462
rect 274504 -3782 274686 -3546
rect 274922 -3782 275104 -3546
rect 274504 -3814 275104 -3782
rect 278204 675694 278804 709082
rect 278204 675458 278386 675694
rect 278622 675458 278804 675694
rect 278204 639694 278804 675458
rect 278204 639458 278386 639694
rect 278622 639458 278804 639694
rect 278204 603694 278804 639458
rect 278204 603458 278386 603694
rect 278622 603458 278804 603694
rect 278204 567694 278804 603458
rect 278204 567458 278386 567694
rect 278622 567458 278804 567694
rect 278204 531694 278804 567458
rect 278204 531458 278386 531694
rect 278622 531458 278804 531694
rect 278204 495694 278804 531458
rect 278204 495458 278386 495694
rect 278622 495458 278804 495694
rect 278204 459694 278804 495458
rect 278204 459458 278386 459694
rect 278622 459458 278804 459694
rect 278204 423694 278804 459458
rect 278204 423458 278386 423694
rect 278622 423458 278804 423694
rect 278204 387694 278804 423458
rect 278204 387458 278386 387694
rect 278622 387458 278804 387694
rect 278204 351694 278804 387458
rect 278204 351458 278386 351694
rect 278622 351458 278804 351694
rect 278204 315694 278804 351458
rect 278204 315458 278386 315694
rect 278622 315458 278804 315694
rect 278204 279694 278804 315458
rect 278204 279458 278386 279694
rect 278622 279458 278804 279694
rect 278204 243694 278804 279458
rect 278204 243458 278386 243694
rect 278622 243458 278804 243694
rect 278204 207694 278804 243458
rect 278204 207458 278386 207694
rect 278622 207458 278804 207694
rect 278204 171694 278804 207458
rect 278204 171458 278386 171694
rect 278622 171458 278804 171694
rect 278204 135694 278804 171458
rect 278204 135458 278386 135694
rect 278622 135458 278804 135694
rect 278204 99694 278804 135458
rect 278204 99458 278386 99694
rect 278622 99458 278804 99694
rect 278204 63694 278804 99458
rect 278204 63458 278386 63694
rect 278622 63458 278804 63694
rect 278204 27694 278804 63458
rect 278204 27458 278386 27694
rect 278622 27458 278804 27694
rect 278204 -5146 278804 27458
rect 278204 -5382 278386 -5146
rect 278622 -5382 278804 -5146
rect 278204 -5466 278804 -5382
rect 278204 -5702 278386 -5466
rect 278622 -5702 278804 -5466
rect 278204 -5734 278804 -5702
rect 281904 679394 282504 711002
rect 299904 710598 300504 711590
rect 299904 710362 300086 710598
rect 300322 710362 300504 710598
rect 299904 710278 300504 710362
rect 299904 710042 300086 710278
rect 300322 710042 300504 710278
rect 296204 708678 296804 709670
rect 296204 708442 296386 708678
rect 296622 708442 296804 708678
rect 296204 708358 296804 708442
rect 296204 708122 296386 708358
rect 296622 708122 296804 708358
rect 292504 706758 293104 707750
rect 292504 706522 292686 706758
rect 292922 706522 293104 706758
rect 292504 706438 293104 706522
rect 292504 706202 292686 706438
rect 292922 706202 293104 706438
rect 281904 679158 282086 679394
rect 282322 679158 282504 679394
rect 281904 643394 282504 679158
rect 281904 643158 282086 643394
rect 282322 643158 282504 643394
rect 281904 607394 282504 643158
rect 281904 607158 282086 607394
rect 282322 607158 282504 607394
rect 281904 571394 282504 607158
rect 281904 571158 282086 571394
rect 282322 571158 282504 571394
rect 281904 535394 282504 571158
rect 281904 535158 282086 535394
rect 282322 535158 282504 535394
rect 281904 499394 282504 535158
rect 281904 499158 282086 499394
rect 282322 499158 282504 499394
rect 281904 463394 282504 499158
rect 281904 463158 282086 463394
rect 282322 463158 282504 463394
rect 281904 427394 282504 463158
rect 281904 427158 282086 427394
rect 282322 427158 282504 427394
rect 281904 391394 282504 427158
rect 281904 391158 282086 391394
rect 282322 391158 282504 391394
rect 281904 355394 282504 391158
rect 281904 355158 282086 355394
rect 282322 355158 282504 355394
rect 281904 319394 282504 355158
rect 281904 319158 282086 319394
rect 282322 319158 282504 319394
rect 281904 283394 282504 319158
rect 281904 283158 282086 283394
rect 282322 283158 282504 283394
rect 281904 247394 282504 283158
rect 281904 247158 282086 247394
rect 282322 247158 282504 247394
rect 281904 211394 282504 247158
rect 281904 211158 282086 211394
rect 282322 211158 282504 211394
rect 281904 175394 282504 211158
rect 281904 175158 282086 175394
rect 282322 175158 282504 175394
rect 281904 139394 282504 175158
rect 281904 139158 282086 139394
rect 282322 139158 282504 139394
rect 281904 103394 282504 139158
rect 281904 103158 282086 103394
rect 282322 103158 282504 103394
rect 281904 67394 282504 103158
rect 281904 67158 282086 67394
rect 282322 67158 282504 67394
rect 281904 31394 282504 67158
rect 281904 31158 282086 31394
rect 282322 31158 282504 31394
rect 263904 -6342 264086 -6106
rect 264322 -6342 264504 -6106
rect 263904 -6426 264504 -6342
rect 263904 -6662 264086 -6426
rect 264322 -6662 264504 -6426
rect 263904 -7654 264504 -6662
rect 281904 -7066 282504 31158
rect 288804 704838 289404 705830
rect 288804 704602 288986 704838
rect 289222 704602 289404 704838
rect 288804 704518 289404 704602
rect 288804 704282 288986 704518
rect 289222 704282 289404 704518
rect 288804 686294 289404 704282
rect 288804 686058 288986 686294
rect 289222 686058 289404 686294
rect 288804 650294 289404 686058
rect 288804 650058 288986 650294
rect 289222 650058 289404 650294
rect 288804 614294 289404 650058
rect 288804 614058 288986 614294
rect 289222 614058 289404 614294
rect 288804 578294 289404 614058
rect 288804 578058 288986 578294
rect 289222 578058 289404 578294
rect 288804 542294 289404 578058
rect 288804 542058 288986 542294
rect 289222 542058 289404 542294
rect 288804 506294 289404 542058
rect 288804 506058 288986 506294
rect 289222 506058 289404 506294
rect 288804 470294 289404 506058
rect 288804 470058 288986 470294
rect 289222 470058 289404 470294
rect 288804 434294 289404 470058
rect 288804 434058 288986 434294
rect 289222 434058 289404 434294
rect 288804 398294 289404 434058
rect 288804 398058 288986 398294
rect 289222 398058 289404 398294
rect 288804 362294 289404 398058
rect 288804 362058 288986 362294
rect 289222 362058 289404 362294
rect 288804 326294 289404 362058
rect 288804 326058 288986 326294
rect 289222 326058 289404 326294
rect 288804 290294 289404 326058
rect 288804 290058 288986 290294
rect 289222 290058 289404 290294
rect 288804 254294 289404 290058
rect 288804 254058 288986 254294
rect 289222 254058 289404 254294
rect 288804 218294 289404 254058
rect 288804 218058 288986 218294
rect 289222 218058 289404 218294
rect 288804 182294 289404 218058
rect 288804 182058 288986 182294
rect 289222 182058 289404 182294
rect 288804 146294 289404 182058
rect 288804 146058 288986 146294
rect 289222 146058 289404 146294
rect 288804 110294 289404 146058
rect 288804 110058 288986 110294
rect 289222 110058 289404 110294
rect 288804 74294 289404 110058
rect 288804 74058 288986 74294
rect 289222 74058 289404 74294
rect 288804 38294 289404 74058
rect 288804 38058 288986 38294
rect 289222 38058 289404 38294
rect 288804 2294 289404 38058
rect 288804 2058 288986 2294
rect 289222 2058 289404 2294
rect 288804 -346 289404 2058
rect 288804 -582 288986 -346
rect 289222 -582 289404 -346
rect 288804 -666 289404 -582
rect 288804 -902 288986 -666
rect 289222 -902 289404 -666
rect 288804 -1894 289404 -902
rect 292504 689994 293104 706202
rect 292504 689758 292686 689994
rect 292922 689758 293104 689994
rect 292504 653994 293104 689758
rect 292504 653758 292686 653994
rect 292922 653758 293104 653994
rect 292504 617994 293104 653758
rect 292504 617758 292686 617994
rect 292922 617758 293104 617994
rect 292504 581994 293104 617758
rect 292504 581758 292686 581994
rect 292922 581758 293104 581994
rect 292504 545994 293104 581758
rect 292504 545758 292686 545994
rect 292922 545758 293104 545994
rect 292504 509994 293104 545758
rect 292504 509758 292686 509994
rect 292922 509758 293104 509994
rect 292504 473994 293104 509758
rect 292504 473758 292686 473994
rect 292922 473758 293104 473994
rect 292504 437994 293104 473758
rect 292504 437758 292686 437994
rect 292922 437758 293104 437994
rect 292504 401994 293104 437758
rect 292504 401758 292686 401994
rect 292922 401758 293104 401994
rect 292504 365994 293104 401758
rect 292504 365758 292686 365994
rect 292922 365758 293104 365994
rect 292504 329994 293104 365758
rect 292504 329758 292686 329994
rect 292922 329758 293104 329994
rect 292504 293994 293104 329758
rect 292504 293758 292686 293994
rect 292922 293758 293104 293994
rect 292504 257994 293104 293758
rect 292504 257758 292686 257994
rect 292922 257758 293104 257994
rect 292504 221994 293104 257758
rect 292504 221758 292686 221994
rect 292922 221758 293104 221994
rect 292504 185994 293104 221758
rect 292504 185758 292686 185994
rect 292922 185758 293104 185994
rect 292504 149994 293104 185758
rect 292504 149758 292686 149994
rect 292922 149758 293104 149994
rect 292504 113994 293104 149758
rect 292504 113758 292686 113994
rect 292922 113758 293104 113994
rect 292504 77994 293104 113758
rect 292504 77758 292686 77994
rect 292922 77758 293104 77994
rect 292504 41994 293104 77758
rect 292504 41758 292686 41994
rect 292922 41758 293104 41994
rect 292504 5994 293104 41758
rect 292504 5758 292686 5994
rect 292922 5758 293104 5994
rect 292504 -2266 293104 5758
rect 292504 -2502 292686 -2266
rect 292922 -2502 293104 -2266
rect 292504 -2586 293104 -2502
rect 292504 -2822 292686 -2586
rect 292922 -2822 293104 -2586
rect 292504 -3814 293104 -2822
rect 296204 693694 296804 708122
rect 296204 693458 296386 693694
rect 296622 693458 296804 693694
rect 296204 657694 296804 693458
rect 296204 657458 296386 657694
rect 296622 657458 296804 657694
rect 296204 621694 296804 657458
rect 296204 621458 296386 621694
rect 296622 621458 296804 621694
rect 296204 585694 296804 621458
rect 296204 585458 296386 585694
rect 296622 585458 296804 585694
rect 296204 549694 296804 585458
rect 296204 549458 296386 549694
rect 296622 549458 296804 549694
rect 296204 513694 296804 549458
rect 296204 513458 296386 513694
rect 296622 513458 296804 513694
rect 296204 477694 296804 513458
rect 296204 477458 296386 477694
rect 296622 477458 296804 477694
rect 296204 441694 296804 477458
rect 296204 441458 296386 441694
rect 296622 441458 296804 441694
rect 296204 405694 296804 441458
rect 296204 405458 296386 405694
rect 296622 405458 296804 405694
rect 296204 369694 296804 405458
rect 296204 369458 296386 369694
rect 296622 369458 296804 369694
rect 296204 333694 296804 369458
rect 296204 333458 296386 333694
rect 296622 333458 296804 333694
rect 296204 297694 296804 333458
rect 296204 297458 296386 297694
rect 296622 297458 296804 297694
rect 296204 261694 296804 297458
rect 296204 261458 296386 261694
rect 296622 261458 296804 261694
rect 296204 225694 296804 261458
rect 296204 225458 296386 225694
rect 296622 225458 296804 225694
rect 296204 189694 296804 225458
rect 296204 189458 296386 189694
rect 296622 189458 296804 189694
rect 296204 153694 296804 189458
rect 296204 153458 296386 153694
rect 296622 153458 296804 153694
rect 296204 117694 296804 153458
rect 296204 117458 296386 117694
rect 296622 117458 296804 117694
rect 296204 81694 296804 117458
rect 296204 81458 296386 81694
rect 296622 81458 296804 81694
rect 296204 45694 296804 81458
rect 296204 45458 296386 45694
rect 296622 45458 296804 45694
rect 296204 9694 296804 45458
rect 296204 9458 296386 9694
rect 296622 9458 296804 9694
rect 296204 -4186 296804 9458
rect 296204 -4422 296386 -4186
rect 296622 -4422 296804 -4186
rect 296204 -4506 296804 -4422
rect 296204 -4742 296386 -4506
rect 296622 -4742 296804 -4506
rect 296204 -5734 296804 -4742
rect 299904 697394 300504 710042
rect 317904 711558 318504 711590
rect 317904 711322 318086 711558
rect 318322 711322 318504 711558
rect 317904 711238 318504 711322
rect 317904 711002 318086 711238
rect 318322 711002 318504 711238
rect 314204 709638 314804 709670
rect 314204 709402 314386 709638
rect 314622 709402 314804 709638
rect 314204 709318 314804 709402
rect 314204 709082 314386 709318
rect 314622 709082 314804 709318
rect 310504 707718 311104 707750
rect 310504 707482 310686 707718
rect 310922 707482 311104 707718
rect 310504 707398 311104 707482
rect 310504 707162 310686 707398
rect 310922 707162 311104 707398
rect 299904 697158 300086 697394
rect 300322 697158 300504 697394
rect 299904 661394 300504 697158
rect 299904 661158 300086 661394
rect 300322 661158 300504 661394
rect 299904 625394 300504 661158
rect 299904 625158 300086 625394
rect 300322 625158 300504 625394
rect 299904 589394 300504 625158
rect 299904 589158 300086 589394
rect 300322 589158 300504 589394
rect 299904 553394 300504 589158
rect 299904 553158 300086 553394
rect 300322 553158 300504 553394
rect 299904 517394 300504 553158
rect 299904 517158 300086 517394
rect 300322 517158 300504 517394
rect 299904 481394 300504 517158
rect 299904 481158 300086 481394
rect 300322 481158 300504 481394
rect 299904 445394 300504 481158
rect 299904 445158 300086 445394
rect 300322 445158 300504 445394
rect 299904 409394 300504 445158
rect 299904 409158 300086 409394
rect 300322 409158 300504 409394
rect 299904 373394 300504 409158
rect 299904 373158 300086 373394
rect 300322 373158 300504 373394
rect 299904 337394 300504 373158
rect 299904 337158 300086 337394
rect 300322 337158 300504 337394
rect 299904 301394 300504 337158
rect 299904 301158 300086 301394
rect 300322 301158 300504 301394
rect 299904 265394 300504 301158
rect 299904 265158 300086 265394
rect 300322 265158 300504 265394
rect 299904 229394 300504 265158
rect 299904 229158 300086 229394
rect 300322 229158 300504 229394
rect 299904 193394 300504 229158
rect 299904 193158 300086 193394
rect 300322 193158 300504 193394
rect 299904 157394 300504 193158
rect 299904 157158 300086 157394
rect 300322 157158 300504 157394
rect 299904 121394 300504 157158
rect 299904 121158 300086 121394
rect 300322 121158 300504 121394
rect 299904 85394 300504 121158
rect 299904 85158 300086 85394
rect 300322 85158 300504 85394
rect 299904 49394 300504 85158
rect 299904 49158 300086 49394
rect 300322 49158 300504 49394
rect 299904 13394 300504 49158
rect 299904 13158 300086 13394
rect 300322 13158 300504 13394
rect 281904 -7302 282086 -7066
rect 282322 -7302 282504 -7066
rect 281904 -7386 282504 -7302
rect 281904 -7622 282086 -7386
rect 282322 -7622 282504 -7386
rect 281904 -7654 282504 -7622
rect 299904 -6106 300504 13158
rect 306804 705798 307404 705830
rect 306804 705562 306986 705798
rect 307222 705562 307404 705798
rect 306804 705478 307404 705562
rect 306804 705242 306986 705478
rect 307222 705242 307404 705478
rect 306804 668294 307404 705242
rect 306804 668058 306986 668294
rect 307222 668058 307404 668294
rect 306804 632294 307404 668058
rect 306804 632058 306986 632294
rect 307222 632058 307404 632294
rect 306804 596294 307404 632058
rect 306804 596058 306986 596294
rect 307222 596058 307404 596294
rect 306804 560294 307404 596058
rect 306804 560058 306986 560294
rect 307222 560058 307404 560294
rect 306804 524294 307404 560058
rect 306804 524058 306986 524294
rect 307222 524058 307404 524294
rect 306804 488294 307404 524058
rect 306804 488058 306986 488294
rect 307222 488058 307404 488294
rect 306804 452294 307404 488058
rect 306804 452058 306986 452294
rect 307222 452058 307404 452294
rect 306804 416294 307404 452058
rect 306804 416058 306986 416294
rect 307222 416058 307404 416294
rect 306804 380294 307404 416058
rect 306804 380058 306986 380294
rect 307222 380058 307404 380294
rect 306804 344294 307404 380058
rect 306804 344058 306986 344294
rect 307222 344058 307404 344294
rect 306804 308294 307404 344058
rect 306804 308058 306986 308294
rect 307222 308058 307404 308294
rect 306804 272294 307404 308058
rect 306804 272058 306986 272294
rect 307222 272058 307404 272294
rect 306804 236294 307404 272058
rect 306804 236058 306986 236294
rect 307222 236058 307404 236294
rect 306804 200294 307404 236058
rect 306804 200058 306986 200294
rect 307222 200058 307404 200294
rect 306804 164294 307404 200058
rect 306804 164058 306986 164294
rect 307222 164058 307404 164294
rect 306804 128294 307404 164058
rect 306804 128058 306986 128294
rect 307222 128058 307404 128294
rect 306804 92294 307404 128058
rect 306804 92058 306986 92294
rect 307222 92058 307404 92294
rect 306804 56294 307404 92058
rect 306804 56058 306986 56294
rect 307222 56058 307404 56294
rect 306804 20294 307404 56058
rect 306804 20058 306986 20294
rect 307222 20058 307404 20294
rect 306804 -1306 307404 20058
rect 306804 -1542 306986 -1306
rect 307222 -1542 307404 -1306
rect 306804 -1626 307404 -1542
rect 306804 -1862 306986 -1626
rect 307222 -1862 307404 -1626
rect 306804 -1894 307404 -1862
rect 310504 671994 311104 707162
rect 310504 671758 310686 671994
rect 310922 671758 311104 671994
rect 310504 635994 311104 671758
rect 310504 635758 310686 635994
rect 310922 635758 311104 635994
rect 310504 599994 311104 635758
rect 310504 599758 310686 599994
rect 310922 599758 311104 599994
rect 310504 563994 311104 599758
rect 310504 563758 310686 563994
rect 310922 563758 311104 563994
rect 310504 527994 311104 563758
rect 310504 527758 310686 527994
rect 310922 527758 311104 527994
rect 310504 491994 311104 527758
rect 310504 491758 310686 491994
rect 310922 491758 311104 491994
rect 310504 455994 311104 491758
rect 310504 455758 310686 455994
rect 310922 455758 311104 455994
rect 310504 419994 311104 455758
rect 310504 419758 310686 419994
rect 310922 419758 311104 419994
rect 310504 383994 311104 419758
rect 310504 383758 310686 383994
rect 310922 383758 311104 383994
rect 310504 347994 311104 383758
rect 310504 347758 310686 347994
rect 310922 347758 311104 347994
rect 310504 311994 311104 347758
rect 310504 311758 310686 311994
rect 310922 311758 311104 311994
rect 310504 275994 311104 311758
rect 310504 275758 310686 275994
rect 310922 275758 311104 275994
rect 310504 239994 311104 275758
rect 310504 239758 310686 239994
rect 310922 239758 311104 239994
rect 310504 203994 311104 239758
rect 310504 203758 310686 203994
rect 310922 203758 311104 203994
rect 310504 167994 311104 203758
rect 310504 167758 310686 167994
rect 310922 167758 311104 167994
rect 310504 131994 311104 167758
rect 310504 131758 310686 131994
rect 310922 131758 311104 131994
rect 310504 95994 311104 131758
rect 310504 95758 310686 95994
rect 310922 95758 311104 95994
rect 310504 59994 311104 95758
rect 310504 59758 310686 59994
rect 310922 59758 311104 59994
rect 310504 23994 311104 59758
rect 310504 23758 310686 23994
rect 310922 23758 311104 23994
rect 310504 -3226 311104 23758
rect 310504 -3462 310686 -3226
rect 310922 -3462 311104 -3226
rect 310504 -3546 311104 -3462
rect 310504 -3782 310686 -3546
rect 310922 -3782 311104 -3546
rect 310504 -3814 311104 -3782
rect 314204 675694 314804 709082
rect 314204 675458 314386 675694
rect 314622 675458 314804 675694
rect 314204 639694 314804 675458
rect 314204 639458 314386 639694
rect 314622 639458 314804 639694
rect 314204 603694 314804 639458
rect 314204 603458 314386 603694
rect 314622 603458 314804 603694
rect 314204 567694 314804 603458
rect 314204 567458 314386 567694
rect 314622 567458 314804 567694
rect 314204 531694 314804 567458
rect 314204 531458 314386 531694
rect 314622 531458 314804 531694
rect 314204 495694 314804 531458
rect 314204 495458 314386 495694
rect 314622 495458 314804 495694
rect 314204 459694 314804 495458
rect 314204 459458 314386 459694
rect 314622 459458 314804 459694
rect 314204 423694 314804 459458
rect 314204 423458 314386 423694
rect 314622 423458 314804 423694
rect 314204 387694 314804 423458
rect 314204 387458 314386 387694
rect 314622 387458 314804 387694
rect 314204 351694 314804 387458
rect 314204 351458 314386 351694
rect 314622 351458 314804 351694
rect 314204 315694 314804 351458
rect 314204 315458 314386 315694
rect 314622 315458 314804 315694
rect 314204 279694 314804 315458
rect 314204 279458 314386 279694
rect 314622 279458 314804 279694
rect 314204 243694 314804 279458
rect 314204 243458 314386 243694
rect 314622 243458 314804 243694
rect 314204 207694 314804 243458
rect 314204 207458 314386 207694
rect 314622 207458 314804 207694
rect 314204 171694 314804 207458
rect 314204 171458 314386 171694
rect 314622 171458 314804 171694
rect 314204 135694 314804 171458
rect 314204 135458 314386 135694
rect 314622 135458 314804 135694
rect 314204 99694 314804 135458
rect 314204 99458 314386 99694
rect 314622 99458 314804 99694
rect 314204 63694 314804 99458
rect 314204 63458 314386 63694
rect 314622 63458 314804 63694
rect 314204 27694 314804 63458
rect 314204 27458 314386 27694
rect 314622 27458 314804 27694
rect 314204 -5146 314804 27458
rect 314204 -5382 314386 -5146
rect 314622 -5382 314804 -5146
rect 314204 -5466 314804 -5382
rect 314204 -5702 314386 -5466
rect 314622 -5702 314804 -5466
rect 314204 -5734 314804 -5702
rect 317904 679394 318504 711002
rect 335904 710598 336504 711590
rect 335904 710362 336086 710598
rect 336322 710362 336504 710598
rect 335904 710278 336504 710362
rect 335904 710042 336086 710278
rect 336322 710042 336504 710278
rect 332204 708678 332804 709670
rect 332204 708442 332386 708678
rect 332622 708442 332804 708678
rect 332204 708358 332804 708442
rect 332204 708122 332386 708358
rect 332622 708122 332804 708358
rect 328504 706758 329104 707750
rect 328504 706522 328686 706758
rect 328922 706522 329104 706758
rect 328504 706438 329104 706522
rect 328504 706202 328686 706438
rect 328922 706202 329104 706438
rect 317904 679158 318086 679394
rect 318322 679158 318504 679394
rect 317904 643394 318504 679158
rect 317904 643158 318086 643394
rect 318322 643158 318504 643394
rect 317904 607394 318504 643158
rect 317904 607158 318086 607394
rect 318322 607158 318504 607394
rect 317904 571394 318504 607158
rect 317904 571158 318086 571394
rect 318322 571158 318504 571394
rect 317904 535394 318504 571158
rect 317904 535158 318086 535394
rect 318322 535158 318504 535394
rect 317904 499394 318504 535158
rect 317904 499158 318086 499394
rect 318322 499158 318504 499394
rect 317904 463394 318504 499158
rect 317904 463158 318086 463394
rect 318322 463158 318504 463394
rect 317904 427394 318504 463158
rect 317904 427158 318086 427394
rect 318322 427158 318504 427394
rect 317904 391394 318504 427158
rect 317904 391158 318086 391394
rect 318322 391158 318504 391394
rect 317904 355394 318504 391158
rect 317904 355158 318086 355394
rect 318322 355158 318504 355394
rect 317904 319394 318504 355158
rect 317904 319158 318086 319394
rect 318322 319158 318504 319394
rect 317904 283394 318504 319158
rect 317904 283158 318086 283394
rect 318322 283158 318504 283394
rect 317904 247394 318504 283158
rect 317904 247158 318086 247394
rect 318322 247158 318504 247394
rect 317904 211394 318504 247158
rect 317904 211158 318086 211394
rect 318322 211158 318504 211394
rect 317904 175394 318504 211158
rect 317904 175158 318086 175394
rect 318322 175158 318504 175394
rect 317904 139394 318504 175158
rect 317904 139158 318086 139394
rect 318322 139158 318504 139394
rect 317904 103394 318504 139158
rect 317904 103158 318086 103394
rect 318322 103158 318504 103394
rect 317904 67394 318504 103158
rect 317904 67158 318086 67394
rect 318322 67158 318504 67394
rect 317904 31394 318504 67158
rect 317904 31158 318086 31394
rect 318322 31158 318504 31394
rect 299904 -6342 300086 -6106
rect 300322 -6342 300504 -6106
rect 299904 -6426 300504 -6342
rect 299904 -6662 300086 -6426
rect 300322 -6662 300504 -6426
rect 299904 -7654 300504 -6662
rect 317904 -7066 318504 31158
rect 324804 704838 325404 705830
rect 324804 704602 324986 704838
rect 325222 704602 325404 704838
rect 324804 704518 325404 704602
rect 324804 704282 324986 704518
rect 325222 704282 325404 704518
rect 324804 686294 325404 704282
rect 324804 686058 324986 686294
rect 325222 686058 325404 686294
rect 324804 650294 325404 686058
rect 324804 650058 324986 650294
rect 325222 650058 325404 650294
rect 324804 614294 325404 650058
rect 324804 614058 324986 614294
rect 325222 614058 325404 614294
rect 324804 578294 325404 614058
rect 324804 578058 324986 578294
rect 325222 578058 325404 578294
rect 324804 542294 325404 578058
rect 324804 542058 324986 542294
rect 325222 542058 325404 542294
rect 324804 506294 325404 542058
rect 324804 506058 324986 506294
rect 325222 506058 325404 506294
rect 324804 470294 325404 506058
rect 324804 470058 324986 470294
rect 325222 470058 325404 470294
rect 324804 434294 325404 470058
rect 324804 434058 324986 434294
rect 325222 434058 325404 434294
rect 324804 398294 325404 434058
rect 324804 398058 324986 398294
rect 325222 398058 325404 398294
rect 324804 362294 325404 398058
rect 324804 362058 324986 362294
rect 325222 362058 325404 362294
rect 324804 326294 325404 362058
rect 324804 326058 324986 326294
rect 325222 326058 325404 326294
rect 324804 290294 325404 326058
rect 324804 290058 324986 290294
rect 325222 290058 325404 290294
rect 324804 254294 325404 290058
rect 324804 254058 324986 254294
rect 325222 254058 325404 254294
rect 324804 218294 325404 254058
rect 324804 218058 324986 218294
rect 325222 218058 325404 218294
rect 324804 182294 325404 218058
rect 324804 182058 324986 182294
rect 325222 182058 325404 182294
rect 324804 146294 325404 182058
rect 324804 146058 324986 146294
rect 325222 146058 325404 146294
rect 324804 110294 325404 146058
rect 324804 110058 324986 110294
rect 325222 110058 325404 110294
rect 324804 74294 325404 110058
rect 324804 74058 324986 74294
rect 325222 74058 325404 74294
rect 324804 38294 325404 74058
rect 324804 38058 324986 38294
rect 325222 38058 325404 38294
rect 324804 2294 325404 38058
rect 324804 2058 324986 2294
rect 325222 2058 325404 2294
rect 324804 -346 325404 2058
rect 324804 -582 324986 -346
rect 325222 -582 325404 -346
rect 324804 -666 325404 -582
rect 324804 -902 324986 -666
rect 325222 -902 325404 -666
rect 324804 -1894 325404 -902
rect 328504 689994 329104 706202
rect 328504 689758 328686 689994
rect 328922 689758 329104 689994
rect 328504 653994 329104 689758
rect 328504 653758 328686 653994
rect 328922 653758 329104 653994
rect 328504 617994 329104 653758
rect 328504 617758 328686 617994
rect 328922 617758 329104 617994
rect 328504 581994 329104 617758
rect 328504 581758 328686 581994
rect 328922 581758 329104 581994
rect 328504 545994 329104 581758
rect 328504 545758 328686 545994
rect 328922 545758 329104 545994
rect 328504 509994 329104 545758
rect 328504 509758 328686 509994
rect 328922 509758 329104 509994
rect 328504 473994 329104 509758
rect 328504 473758 328686 473994
rect 328922 473758 329104 473994
rect 328504 437994 329104 473758
rect 328504 437758 328686 437994
rect 328922 437758 329104 437994
rect 328504 401994 329104 437758
rect 328504 401758 328686 401994
rect 328922 401758 329104 401994
rect 328504 365994 329104 401758
rect 328504 365758 328686 365994
rect 328922 365758 329104 365994
rect 328504 329994 329104 365758
rect 328504 329758 328686 329994
rect 328922 329758 329104 329994
rect 328504 293994 329104 329758
rect 328504 293758 328686 293994
rect 328922 293758 329104 293994
rect 328504 257994 329104 293758
rect 328504 257758 328686 257994
rect 328922 257758 329104 257994
rect 328504 221994 329104 257758
rect 328504 221758 328686 221994
rect 328922 221758 329104 221994
rect 328504 185994 329104 221758
rect 328504 185758 328686 185994
rect 328922 185758 329104 185994
rect 328504 149994 329104 185758
rect 328504 149758 328686 149994
rect 328922 149758 329104 149994
rect 328504 113994 329104 149758
rect 328504 113758 328686 113994
rect 328922 113758 329104 113994
rect 328504 77994 329104 113758
rect 328504 77758 328686 77994
rect 328922 77758 329104 77994
rect 328504 41994 329104 77758
rect 328504 41758 328686 41994
rect 328922 41758 329104 41994
rect 328504 5994 329104 41758
rect 328504 5758 328686 5994
rect 328922 5758 329104 5994
rect 328504 -2266 329104 5758
rect 328504 -2502 328686 -2266
rect 328922 -2502 329104 -2266
rect 328504 -2586 329104 -2502
rect 328504 -2822 328686 -2586
rect 328922 -2822 329104 -2586
rect 328504 -3814 329104 -2822
rect 332204 693694 332804 708122
rect 332204 693458 332386 693694
rect 332622 693458 332804 693694
rect 332204 657694 332804 693458
rect 332204 657458 332386 657694
rect 332622 657458 332804 657694
rect 332204 621694 332804 657458
rect 332204 621458 332386 621694
rect 332622 621458 332804 621694
rect 332204 585694 332804 621458
rect 332204 585458 332386 585694
rect 332622 585458 332804 585694
rect 332204 549694 332804 585458
rect 332204 549458 332386 549694
rect 332622 549458 332804 549694
rect 332204 513694 332804 549458
rect 332204 513458 332386 513694
rect 332622 513458 332804 513694
rect 332204 477694 332804 513458
rect 332204 477458 332386 477694
rect 332622 477458 332804 477694
rect 332204 441694 332804 477458
rect 332204 441458 332386 441694
rect 332622 441458 332804 441694
rect 332204 405694 332804 441458
rect 332204 405458 332386 405694
rect 332622 405458 332804 405694
rect 332204 369694 332804 405458
rect 332204 369458 332386 369694
rect 332622 369458 332804 369694
rect 332204 333694 332804 369458
rect 332204 333458 332386 333694
rect 332622 333458 332804 333694
rect 332204 297694 332804 333458
rect 332204 297458 332386 297694
rect 332622 297458 332804 297694
rect 332204 261694 332804 297458
rect 332204 261458 332386 261694
rect 332622 261458 332804 261694
rect 332204 225694 332804 261458
rect 332204 225458 332386 225694
rect 332622 225458 332804 225694
rect 332204 189694 332804 225458
rect 332204 189458 332386 189694
rect 332622 189458 332804 189694
rect 332204 153694 332804 189458
rect 332204 153458 332386 153694
rect 332622 153458 332804 153694
rect 332204 117694 332804 153458
rect 332204 117458 332386 117694
rect 332622 117458 332804 117694
rect 332204 81694 332804 117458
rect 332204 81458 332386 81694
rect 332622 81458 332804 81694
rect 332204 45694 332804 81458
rect 332204 45458 332386 45694
rect 332622 45458 332804 45694
rect 332204 9694 332804 45458
rect 332204 9458 332386 9694
rect 332622 9458 332804 9694
rect 332204 -4186 332804 9458
rect 332204 -4422 332386 -4186
rect 332622 -4422 332804 -4186
rect 332204 -4506 332804 -4422
rect 332204 -4742 332386 -4506
rect 332622 -4742 332804 -4506
rect 332204 -5734 332804 -4742
rect 335904 697394 336504 710042
rect 353904 711558 354504 711590
rect 353904 711322 354086 711558
rect 354322 711322 354504 711558
rect 353904 711238 354504 711322
rect 353904 711002 354086 711238
rect 354322 711002 354504 711238
rect 350204 709638 350804 709670
rect 350204 709402 350386 709638
rect 350622 709402 350804 709638
rect 350204 709318 350804 709402
rect 350204 709082 350386 709318
rect 350622 709082 350804 709318
rect 346504 707718 347104 707750
rect 346504 707482 346686 707718
rect 346922 707482 347104 707718
rect 346504 707398 347104 707482
rect 346504 707162 346686 707398
rect 346922 707162 347104 707398
rect 335904 697158 336086 697394
rect 336322 697158 336504 697394
rect 335904 661394 336504 697158
rect 335904 661158 336086 661394
rect 336322 661158 336504 661394
rect 335904 625394 336504 661158
rect 335904 625158 336086 625394
rect 336322 625158 336504 625394
rect 335904 589394 336504 625158
rect 335904 589158 336086 589394
rect 336322 589158 336504 589394
rect 335904 553394 336504 589158
rect 335904 553158 336086 553394
rect 336322 553158 336504 553394
rect 335904 517394 336504 553158
rect 335904 517158 336086 517394
rect 336322 517158 336504 517394
rect 335904 481394 336504 517158
rect 335904 481158 336086 481394
rect 336322 481158 336504 481394
rect 335904 445394 336504 481158
rect 335904 445158 336086 445394
rect 336322 445158 336504 445394
rect 335904 409394 336504 445158
rect 342804 705798 343404 705830
rect 342804 705562 342986 705798
rect 343222 705562 343404 705798
rect 342804 705478 343404 705562
rect 342804 705242 342986 705478
rect 343222 705242 343404 705478
rect 342804 668294 343404 705242
rect 342804 668058 342986 668294
rect 343222 668058 343404 668294
rect 342804 632294 343404 668058
rect 342804 632058 342986 632294
rect 343222 632058 343404 632294
rect 342804 596294 343404 632058
rect 342804 596058 342986 596294
rect 343222 596058 343404 596294
rect 342804 560294 343404 596058
rect 342804 560058 342986 560294
rect 343222 560058 343404 560294
rect 342804 524294 343404 560058
rect 342804 524058 342986 524294
rect 343222 524058 343404 524294
rect 342804 488294 343404 524058
rect 342804 488058 342986 488294
rect 343222 488058 343404 488294
rect 342804 452294 343404 488058
rect 342804 452058 342986 452294
rect 343222 452058 343404 452294
rect 342804 425308 343404 452058
rect 346504 671994 347104 707162
rect 346504 671758 346686 671994
rect 346922 671758 347104 671994
rect 346504 635994 347104 671758
rect 346504 635758 346686 635994
rect 346922 635758 347104 635994
rect 346504 599994 347104 635758
rect 346504 599758 346686 599994
rect 346922 599758 347104 599994
rect 346504 563994 347104 599758
rect 346504 563758 346686 563994
rect 346922 563758 347104 563994
rect 346504 527994 347104 563758
rect 346504 527758 346686 527994
rect 346922 527758 347104 527994
rect 346504 491994 347104 527758
rect 346504 491758 346686 491994
rect 346922 491758 347104 491994
rect 346504 455994 347104 491758
rect 346504 455758 346686 455994
rect 346922 455758 347104 455994
rect 346504 425308 347104 455758
rect 350204 675694 350804 709082
rect 350204 675458 350386 675694
rect 350622 675458 350804 675694
rect 350204 639694 350804 675458
rect 350204 639458 350386 639694
rect 350622 639458 350804 639694
rect 350204 603694 350804 639458
rect 350204 603458 350386 603694
rect 350622 603458 350804 603694
rect 350204 567694 350804 603458
rect 350204 567458 350386 567694
rect 350622 567458 350804 567694
rect 350204 531694 350804 567458
rect 350204 531458 350386 531694
rect 350622 531458 350804 531694
rect 350204 495694 350804 531458
rect 350204 495458 350386 495694
rect 350622 495458 350804 495694
rect 350204 459694 350804 495458
rect 350204 459458 350386 459694
rect 350622 459458 350804 459694
rect 350204 425308 350804 459458
rect 353904 679394 354504 711002
rect 371904 710598 372504 711590
rect 371904 710362 372086 710598
rect 372322 710362 372504 710598
rect 371904 710278 372504 710362
rect 371904 710042 372086 710278
rect 372322 710042 372504 710278
rect 368204 708678 368804 709670
rect 368204 708442 368386 708678
rect 368622 708442 368804 708678
rect 368204 708358 368804 708442
rect 368204 708122 368386 708358
rect 368622 708122 368804 708358
rect 364504 706758 365104 707750
rect 364504 706522 364686 706758
rect 364922 706522 365104 706758
rect 364504 706438 365104 706522
rect 364504 706202 364686 706438
rect 364922 706202 365104 706438
rect 353904 679158 354086 679394
rect 354322 679158 354504 679394
rect 353904 643394 354504 679158
rect 353904 643158 354086 643394
rect 354322 643158 354504 643394
rect 353904 607394 354504 643158
rect 353904 607158 354086 607394
rect 354322 607158 354504 607394
rect 353904 571394 354504 607158
rect 353904 571158 354086 571394
rect 354322 571158 354504 571394
rect 353904 535394 354504 571158
rect 353904 535158 354086 535394
rect 354322 535158 354504 535394
rect 353904 499394 354504 535158
rect 353904 499158 354086 499394
rect 354322 499158 354504 499394
rect 353904 463394 354504 499158
rect 353904 463158 354086 463394
rect 354322 463158 354504 463394
rect 353904 427394 354504 463158
rect 353904 427158 354086 427394
rect 354322 427158 354504 427394
rect 353904 425308 354504 427158
rect 360804 704838 361404 705830
rect 360804 704602 360986 704838
rect 361222 704602 361404 704838
rect 360804 704518 361404 704602
rect 360804 704282 360986 704518
rect 361222 704282 361404 704518
rect 360804 686294 361404 704282
rect 360804 686058 360986 686294
rect 361222 686058 361404 686294
rect 360804 650294 361404 686058
rect 360804 650058 360986 650294
rect 361222 650058 361404 650294
rect 360804 614294 361404 650058
rect 360804 614058 360986 614294
rect 361222 614058 361404 614294
rect 360804 578294 361404 614058
rect 360804 578058 360986 578294
rect 361222 578058 361404 578294
rect 360804 542294 361404 578058
rect 360804 542058 360986 542294
rect 361222 542058 361404 542294
rect 360804 506294 361404 542058
rect 360804 506058 360986 506294
rect 361222 506058 361404 506294
rect 360804 470294 361404 506058
rect 360804 470058 360986 470294
rect 361222 470058 361404 470294
rect 360804 434294 361404 470058
rect 360804 434058 360986 434294
rect 361222 434058 361404 434294
rect 360804 425308 361404 434058
rect 364504 689994 365104 706202
rect 364504 689758 364686 689994
rect 364922 689758 365104 689994
rect 364504 653994 365104 689758
rect 364504 653758 364686 653994
rect 364922 653758 365104 653994
rect 364504 617994 365104 653758
rect 364504 617758 364686 617994
rect 364922 617758 365104 617994
rect 364504 581994 365104 617758
rect 364504 581758 364686 581994
rect 364922 581758 365104 581994
rect 364504 545994 365104 581758
rect 364504 545758 364686 545994
rect 364922 545758 365104 545994
rect 364504 509994 365104 545758
rect 364504 509758 364686 509994
rect 364922 509758 365104 509994
rect 364504 473994 365104 509758
rect 364504 473758 364686 473994
rect 364922 473758 365104 473994
rect 364504 437994 365104 473758
rect 364504 437758 364686 437994
rect 364922 437758 365104 437994
rect 364504 425308 365104 437758
rect 368204 693694 368804 708122
rect 368204 693458 368386 693694
rect 368622 693458 368804 693694
rect 368204 657694 368804 693458
rect 368204 657458 368386 657694
rect 368622 657458 368804 657694
rect 368204 621694 368804 657458
rect 368204 621458 368386 621694
rect 368622 621458 368804 621694
rect 368204 585694 368804 621458
rect 368204 585458 368386 585694
rect 368622 585458 368804 585694
rect 368204 549694 368804 585458
rect 368204 549458 368386 549694
rect 368622 549458 368804 549694
rect 368204 513694 368804 549458
rect 368204 513458 368386 513694
rect 368622 513458 368804 513694
rect 368204 477694 368804 513458
rect 368204 477458 368386 477694
rect 368622 477458 368804 477694
rect 368204 441694 368804 477458
rect 368204 441458 368386 441694
rect 368622 441458 368804 441694
rect 368204 425308 368804 441458
rect 371904 697394 372504 710042
rect 389904 711558 390504 711590
rect 389904 711322 390086 711558
rect 390322 711322 390504 711558
rect 389904 711238 390504 711322
rect 389904 711002 390086 711238
rect 390322 711002 390504 711238
rect 386204 709638 386804 709670
rect 386204 709402 386386 709638
rect 386622 709402 386804 709638
rect 386204 709318 386804 709402
rect 386204 709082 386386 709318
rect 386622 709082 386804 709318
rect 382504 707718 383104 707750
rect 382504 707482 382686 707718
rect 382922 707482 383104 707718
rect 382504 707398 383104 707482
rect 382504 707162 382686 707398
rect 382922 707162 383104 707398
rect 371904 697158 372086 697394
rect 372322 697158 372504 697394
rect 371904 661394 372504 697158
rect 371904 661158 372086 661394
rect 372322 661158 372504 661394
rect 371904 625394 372504 661158
rect 371904 625158 372086 625394
rect 372322 625158 372504 625394
rect 371904 589394 372504 625158
rect 371904 589158 372086 589394
rect 372322 589158 372504 589394
rect 371904 553394 372504 589158
rect 371904 553158 372086 553394
rect 372322 553158 372504 553394
rect 371904 517394 372504 553158
rect 371904 517158 372086 517394
rect 372322 517158 372504 517394
rect 371904 481394 372504 517158
rect 371904 481158 372086 481394
rect 372322 481158 372504 481394
rect 371904 445394 372504 481158
rect 371904 445158 372086 445394
rect 372322 445158 372504 445394
rect 371904 425308 372504 445158
rect 378804 705798 379404 705830
rect 378804 705562 378986 705798
rect 379222 705562 379404 705798
rect 378804 705478 379404 705562
rect 378804 705242 378986 705478
rect 379222 705242 379404 705478
rect 378804 668294 379404 705242
rect 378804 668058 378986 668294
rect 379222 668058 379404 668294
rect 378804 632294 379404 668058
rect 378804 632058 378986 632294
rect 379222 632058 379404 632294
rect 378804 596294 379404 632058
rect 378804 596058 378986 596294
rect 379222 596058 379404 596294
rect 378804 560294 379404 596058
rect 378804 560058 378986 560294
rect 379222 560058 379404 560294
rect 378804 524294 379404 560058
rect 378804 524058 378986 524294
rect 379222 524058 379404 524294
rect 378804 488294 379404 524058
rect 378804 488058 378986 488294
rect 379222 488058 379404 488294
rect 378804 452294 379404 488058
rect 378804 452058 378986 452294
rect 379222 452058 379404 452294
rect 378804 425308 379404 452058
rect 382504 671994 383104 707162
rect 382504 671758 382686 671994
rect 382922 671758 383104 671994
rect 382504 635994 383104 671758
rect 382504 635758 382686 635994
rect 382922 635758 383104 635994
rect 382504 599994 383104 635758
rect 382504 599758 382686 599994
rect 382922 599758 383104 599994
rect 382504 563994 383104 599758
rect 382504 563758 382686 563994
rect 382922 563758 383104 563994
rect 382504 527994 383104 563758
rect 382504 527758 382686 527994
rect 382922 527758 383104 527994
rect 382504 491994 383104 527758
rect 382504 491758 382686 491994
rect 382922 491758 383104 491994
rect 382504 455994 383104 491758
rect 382504 455758 382686 455994
rect 382922 455758 383104 455994
rect 382504 425308 383104 455758
rect 386204 675694 386804 709082
rect 386204 675458 386386 675694
rect 386622 675458 386804 675694
rect 386204 639694 386804 675458
rect 386204 639458 386386 639694
rect 386622 639458 386804 639694
rect 386204 603694 386804 639458
rect 386204 603458 386386 603694
rect 386622 603458 386804 603694
rect 386204 567694 386804 603458
rect 386204 567458 386386 567694
rect 386622 567458 386804 567694
rect 386204 531694 386804 567458
rect 386204 531458 386386 531694
rect 386622 531458 386804 531694
rect 386204 495694 386804 531458
rect 386204 495458 386386 495694
rect 386622 495458 386804 495694
rect 386204 459694 386804 495458
rect 386204 459458 386386 459694
rect 386622 459458 386804 459694
rect 386204 425308 386804 459458
rect 389904 679394 390504 711002
rect 407904 710598 408504 711590
rect 407904 710362 408086 710598
rect 408322 710362 408504 710598
rect 407904 710278 408504 710362
rect 407904 710042 408086 710278
rect 408322 710042 408504 710278
rect 404204 708678 404804 709670
rect 404204 708442 404386 708678
rect 404622 708442 404804 708678
rect 404204 708358 404804 708442
rect 404204 708122 404386 708358
rect 404622 708122 404804 708358
rect 400504 706758 401104 707750
rect 400504 706522 400686 706758
rect 400922 706522 401104 706758
rect 400504 706438 401104 706522
rect 400504 706202 400686 706438
rect 400922 706202 401104 706438
rect 389904 679158 390086 679394
rect 390322 679158 390504 679394
rect 389904 643394 390504 679158
rect 389904 643158 390086 643394
rect 390322 643158 390504 643394
rect 389904 607394 390504 643158
rect 389904 607158 390086 607394
rect 390322 607158 390504 607394
rect 389904 571394 390504 607158
rect 389904 571158 390086 571394
rect 390322 571158 390504 571394
rect 389904 535394 390504 571158
rect 389904 535158 390086 535394
rect 390322 535158 390504 535394
rect 389904 499394 390504 535158
rect 389904 499158 390086 499394
rect 390322 499158 390504 499394
rect 389904 463394 390504 499158
rect 389904 463158 390086 463394
rect 390322 463158 390504 463394
rect 389904 427394 390504 463158
rect 389904 427158 390086 427394
rect 390322 427158 390504 427394
rect 389904 425308 390504 427158
rect 396804 704838 397404 705830
rect 396804 704602 396986 704838
rect 397222 704602 397404 704838
rect 396804 704518 397404 704602
rect 396804 704282 396986 704518
rect 397222 704282 397404 704518
rect 396804 686294 397404 704282
rect 396804 686058 396986 686294
rect 397222 686058 397404 686294
rect 396804 650294 397404 686058
rect 396804 650058 396986 650294
rect 397222 650058 397404 650294
rect 396804 614294 397404 650058
rect 396804 614058 396986 614294
rect 397222 614058 397404 614294
rect 396804 578294 397404 614058
rect 396804 578058 396986 578294
rect 397222 578058 397404 578294
rect 396804 542294 397404 578058
rect 396804 542058 396986 542294
rect 397222 542058 397404 542294
rect 396804 506294 397404 542058
rect 396804 506058 396986 506294
rect 397222 506058 397404 506294
rect 396804 470294 397404 506058
rect 396804 470058 396986 470294
rect 397222 470058 397404 470294
rect 396804 434294 397404 470058
rect 396804 434058 396986 434294
rect 397222 434058 397404 434294
rect 396804 425308 397404 434058
rect 400504 689994 401104 706202
rect 400504 689758 400686 689994
rect 400922 689758 401104 689994
rect 400504 653994 401104 689758
rect 400504 653758 400686 653994
rect 400922 653758 401104 653994
rect 400504 617994 401104 653758
rect 400504 617758 400686 617994
rect 400922 617758 401104 617994
rect 400504 581994 401104 617758
rect 400504 581758 400686 581994
rect 400922 581758 401104 581994
rect 400504 545994 401104 581758
rect 400504 545758 400686 545994
rect 400922 545758 401104 545994
rect 400504 509994 401104 545758
rect 400504 509758 400686 509994
rect 400922 509758 401104 509994
rect 400504 473994 401104 509758
rect 400504 473758 400686 473994
rect 400922 473758 401104 473994
rect 400504 437994 401104 473758
rect 400504 437758 400686 437994
rect 400922 437758 401104 437994
rect 400504 425308 401104 437758
rect 404204 693694 404804 708122
rect 404204 693458 404386 693694
rect 404622 693458 404804 693694
rect 404204 657694 404804 693458
rect 404204 657458 404386 657694
rect 404622 657458 404804 657694
rect 404204 621694 404804 657458
rect 404204 621458 404386 621694
rect 404622 621458 404804 621694
rect 404204 585694 404804 621458
rect 404204 585458 404386 585694
rect 404622 585458 404804 585694
rect 404204 549694 404804 585458
rect 404204 549458 404386 549694
rect 404622 549458 404804 549694
rect 404204 513694 404804 549458
rect 404204 513458 404386 513694
rect 404622 513458 404804 513694
rect 404204 477694 404804 513458
rect 404204 477458 404386 477694
rect 404622 477458 404804 477694
rect 404204 441694 404804 477458
rect 404204 441458 404386 441694
rect 404622 441458 404804 441694
rect 404204 425308 404804 441458
rect 407904 697394 408504 710042
rect 425904 711558 426504 711590
rect 425904 711322 426086 711558
rect 426322 711322 426504 711558
rect 425904 711238 426504 711322
rect 425904 711002 426086 711238
rect 426322 711002 426504 711238
rect 422204 709638 422804 709670
rect 422204 709402 422386 709638
rect 422622 709402 422804 709638
rect 422204 709318 422804 709402
rect 422204 709082 422386 709318
rect 422622 709082 422804 709318
rect 418504 707718 419104 707750
rect 418504 707482 418686 707718
rect 418922 707482 419104 707718
rect 418504 707398 419104 707482
rect 418504 707162 418686 707398
rect 418922 707162 419104 707398
rect 407904 697158 408086 697394
rect 408322 697158 408504 697394
rect 407904 661394 408504 697158
rect 407904 661158 408086 661394
rect 408322 661158 408504 661394
rect 407904 625394 408504 661158
rect 407904 625158 408086 625394
rect 408322 625158 408504 625394
rect 407904 589394 408504 625158
rect 407904 589158 408086 589394
rect 408322 589158 408504 589394
rect 407904 553394 408504 589158
rect 407904 553158 408086 553394
rect 408322 553158 408504 553394
rect 407904 517394 408504 553158
rect 407904 517158 408086 517394
rect 408322 517158 408504 517394
rect 407904 481394 408504 517158
rect 407904 481158 408086 481394
rect 408322 481158 408504 481394
rect 407904 445394 408504 481158
rect 407904 445158 408086 445394
rect 408322 445158 408504 445394
rect 407904 425308 408504 445158
rect 414804 705798 415404 705830
rect 414804 705562 414986 705798
rect 415222 705562 415404 705798
rect 414804 705478 415404 705562
rect 414804 705242 414986 705478
rect 415222 705242 415404 705478
rect 414804 668294 415404 705242
rect 414804 668058 414986 668294
rect 415222 668058 415404 668294
rect 414804 632294 415404 668058
rect 414804 632058 414986 632294
rect 415222 632058 415404 632294
rect 414804 596294 415404 632058
rect 414804 596058 414986 596294
rect 415222 596058 415404 596294
rect 414804 560294 415404 596058
rect 414804 560058 414986 560294
rect 415222 560058 415404 560294
rect 414804 524294 415404 560058
rect 414804 524058 414986 524294
rect 415222 524058 415404 524294
rect 414804 488294 415404 524058
rect 414804 488058 414986 488294
rect 415222 488058 415404 488294
rect 414804 452294 415404 488058
rect 414804 452058 414986 452294
rect 415222 452058 415404 452294
rect 414804 425308 415404 452058
rect 418504 671994 419104 707162
rect 418504 671758 418686 671994
rect 418922 671758 419104 671994
rect 418504 635994 419104 671758
rect 418504 635758 418686 635994
rect 418922 635758 419104 635994
rect 418504 599994 419104 635758
rect 418504 599758 418686 599994
rect 418922 599758 419104 599994
rect 418504 563994 419104 599758
rect 418504 563758 418686 563994
rect 418922 563758 419104 563994
rect 418504 527994 419104 563758
rect 418504 527758 418686 527994
rect 418922 527758 419104 527994
rect 418504 491994 419104 527758
rect 418504 491758 418686 491994
rect 418922 491758 419104 491994
rect 418504 455994 419104 491758
rect 418504 455758 418686 455994
rect 418922 455758 419104 455994
rect 418504 425308 419104 455758
rect 422204 675694 422804 709082
rect 422204 675458 422386 675694
rect 422622 675458 422804 675694
rect 422204 639694 422804 675458
rect 422204 639458 422386 639694
rect 422622 639458 422804 639694
rect 422204 603694 422804 639458
rect 422204 603458 422386 603694
rect 422622 603458 422804 603694
rect 422204 567694 422804 603458
rect 422204 567458 422386 567694
rect 422622 567458 422804 567694
rect 422204 531694 422804 567458
rect 422204 531458 422386 531694
rect 422622 531458 422804 531694
rect 422204 495694 422804 531458
rect 422204 495458 422386 495694
rect 422622 495458 422804 495694
rect 422204 459694 422804 495458
rect 422204 459458 422386 459694
rect 422622 459458 422804 459694
rect 422204 425308 422804 459458
rect 425904 679394 426504 711002
rect 443904 710598 444504 711590
rect 443904 710362 444086 710598
rect 444322 710362 444504 710598
rect 443904 710278 444504 710362
rect 443904 710042 444086 710278
rect 444322 710042 444504 710278
rect 440204 708678 440804 709670
rect 440204 708442 440386 708678
rect 440622 708442 440804 708678
rect 440204 708358 440804 708442
rect 440204 708122 440386 708358
rect 440622 708122 440804 708358
rect 436504 706758 437104 707750
rect 436504 706522 436686 706758
rect 436922 706522 437104 706758
rect 436504 706438 437104 706522
rect 436504 706202 436686 706438
rect 436922 706202 437104 706438
rect 425904 679158 426086 679394
rect 426322 679158 426504 679394
rect 425904 643394 426504 679158
rect 425904 643158 426086 643394
rect 426322 643158 426504 643394
rect 425904 607394 426504 643158
rect 425904 607158 426086 607394
rect 426322 607158 426504 607394
rect 425904 571394 426504 607158
rect 425904 571158 426086 571394
rect 426322 571158 426504 571394
rect 425904 535394 426504 571158
rect 425904 535158 426086 535394
rect 426322 535158 426504 535394
rect 425904 499394 426504 535158
rect 425904 499158 426086 499394
rect 426322 499158 426504 499394
rect 425904 463394 426504 499158
rect 425904 463158 426086 463394
rect 426322 463158 426504 463394
rect 425904 427394 426504 463158
rect 425904 427158 426086 427394
rect 426322 427158 426504 427394
rect 425904 425308 426504 427158
rect 432804 704838 433404 705830
rect 432804 704602 432986 704838
rect 433222 704602 433404 704838
rect 432804 704518 433404 704602
rect 432804 704282 432986 704518
rect 433222 704282 433404 704518
rect 432804 686294 433404 704282
rect 432804 686058 432986 686294
rect 433222 686058 433404 686294
rect 432804 650294 433404 686058
rect 432804 650058 432986 650294
rect 433222 650058 433404 650294
rect 432804 614294 433404 650058
rect 432804 614058 432986 614294
rect 433222 614058 433404 614294
rect 432804 578294 433404 614058
rect 432804 578058 432986 578294
rect 433222 578058 433404 578294
rect 432804 542294 433404 578058
rect 432804 542058 432986 542294
rect 433222 542058 433404 542294
rect 432804 506294 433404 542058
rect 432804 506058 432986 506294
rect 433222 506058 433404 506294
rect 432804 470294 433404 506058
rect 432804 470058 432986 470294
rect 433222 470058 433404 470294
rect 432804 434294 433404 470058
rect 432804 434058 432986 434294
rect 433222 434058 433404 434294
rect 432804 425308 433404 434058
rect 436504 689994 437104 706202
rect 436504 689758 436686 689994
rect 436922 689758 437104 689994
rect 436504 653994 437104 689758
rect 436504 653758 436686 653994
rect 436922 653758 437104 653994
rect 436504 617994 437104 653758
rect 436504 617758 436686 617994
rect 436922 617758 437104 617994
rect 436504 581994 437104 617758
rect 436504 581758 436686 581994
rect 436922 581758 437104 581994
rect 436504 545994 437104 581758
rect 436504 545758 436686 545994
rect 436922 545758 437104 545994
rect 436504 509994 437104 545758
rect 436504 509758 436686 509994
rect 436922 509758 437104 509994
rect 436504 473994 437104 509758
rect 436504 473758 436686 473994
rect 436922 473758 437104 473994
rect 436504 437994 437104 473758
rect 436504 437758 436686 437994
rect 436922 437758 437104 437994
rect 436504 425308 437104 437758
rect 440204 693694 440804 708122
rect 440204 693458 440386 693694
rect 440622 693458 440804 693694
rect 440204 657694 440804 693458
rect 440204 657458 440386 657694
rect 440622 657458 440804 657694
rect 440204 621694 440804 657458
rect 440204 621458 440386 621694
rect 440622 621458 440804 621694
rect 440204 585694 440804 621458
rect 440204 585458 440386 585694
rect 440622 585458 440804 585694
rect 440204 549694 440804 585458
rect 440204 549458 440386 549694
rect 440622 549458 440804 549694
rect 440204 513694 440804 549458
rect 440204 513458 440386 513694
rect 440622 513458 440804 513694
rect 440204 477694 440804 513458
rect 440204 477458 440386 477694
rect 440622 477458 440804 477694
rect 440204 441694 440804 477458
rect 440204 441458 440386 441694
rect 440622 441458 440804 441694
rect 440204 425308 440804 441458
rect 443904 697394 444504 710042
rect 461904 711558 462504 711590
rect 461904 711322 462086 711558
rect 462322 711322 462504 711558
rect 461904 711238 462504 711322
rect 461904 711002 462086 711238
rect 462322 711002 462504 711238
rect 458204 709638 458804 709670
rect 458204 709402 458386 709638
rect 458622 709402 458804 709638
rect 458204 709318 458804 709402
rect 458204 709082 458386 709318
rect 458622 709082 458804 709318
rect 454504 707718 455104 707750
rect 454504 707482 454686 707718
rect 454922 707482 455104 707718
rect 454504 707398 455104 707482
rect 454504 707162 454686 707398
rect 454922 707162 455104 707398
rect 443904 697158 444086 697394
rect 444322 697158 444504 697394
rect 443904 661394 444504 697158
rect 443904 661158 444086 661394
rect 444322 661158 444504 661394
rect 443904 625394 444504 661158
rect 443904 625158 444086 625394
rect 444322 625158 444504 625394
rect 443904 589394 444504 625158
rect 443904 589158 444086 589394
rect 444322 589158 444504 589394
rect 443904 553394 444504 589158
rect 443904 553158 444086 553394
rect 444322 553158 444504 553394
rect 443904 517394 444504 553158
rect 443904 517158 444086 517394
rect 444322 517158 444504 517394
rect 443904 481394 444504 517158
rect 443904 481158 444086 481394
rect 444322 481158 444504 481394
rect 443904 445394 444504 481158
rect 443904 445158 444086 445394
rect 444322 445158 444504 445394
rect 443904 425308 444504 445158
rect 450804 705798 451404 705830
rect 450804 705562 450986 705798
rect 451222 705562 451404 705798
rect 450804 705478 451404 705562
rect 450804 705242 450986 705478
rect 451222 705242 451404 705478
rect 450804 668294 451404 705242
rect 450804 668058 450986 668294
rect 451222 668058 451404 668294
rect 450804 632294 451404 668058
rect 450804 632058 450986 632294
rect 451222 632058 451404 632294
rect 450804 596294 451404 632058
rect 450804 596058 450986 596294
rect 451222 596058 451404 596294
rect 450804 560294 451404 596058
rect 450804 560058 450986 560294
rect 451222 560058 451404 560294
rect 450804 524294 451404 560058
rect 450804 524058 450986 524294
rect 451222 524058 451404 524294
rect 450804 488294 451404 524058
rect 450804 488058 450986 488294
rect 451222 488058 451404 488294
rect 450804 452294 451404 488058
rect 450804 452058 450986 452294
rect 451222 452058 451404 452294
rect 450804 425308 451404 452058
rect 454504 671994 455104 707162
rect 454504 671758 454686 671994
rect 454922 671758 455104 671994
rect 454504 635994 455104 671758
rect 454504 635758 454686 635994
rect 454922 635758 455104 635994
rect 454504 599994 455104 635758
rect 454504 599758 454686 599994
rect 454922 599758 455104 599994
rect 454504 563994 455104 599758
rect 454504 563758 454686 563994
rect 454922 563758 455104 563994
rect 454504 527994 455104 563758
rect 454504 527758 454686 527994
rect 454922 527758 455104 527994
rect 454504 491994 455104 527758
rect 454504 491758 454686 491994
rect 454922 491758 455104 491994
rect 454504 455994 455104 491758
rect 454504 455758 454686 455994
rect 454922 455758 455104 455994
rect 454504 425308 455104 455758
rect 458204 675694 458804 709082
rect 458204 675458 458386 675694
rect 458622 675458 458804 675694
rect 458204 639694 458804 675458
rect 458204 639458 458386 639694
rect 458622 639458 458804 639694
rect 458204 603694 458804 639458
rect 458204 603458 458386 603694
rect 458622 603458 458804 603694
rect 458204 567694 458804 603458
rect 458204 567458 458386 567694
rect 458622 567458 458804 567694
rect 458204 531694 458804 567458
rect 458204 531458 458386 531694
rect 458622 531458 458804 531694
rect 458204 495694 458804 531458
rect 458204 495458 458386 495694
rect 458622 495458 458804 495694
rect 458204 459694 458804 495458
rect 458204 459458 458386 459694
rect 458622 459458 458804 459694
rect 458204 425308 458804 459458
rect 461904 679394 462504 711002
rect 479904 710598 480504 711590
rect 479904 710362 480086 710598
rect 480322 710362 480504 710598
rect 479904 710278 480504 710362
rect 479904 710042 480086 710278
rect 480322 710042 480504 710278
rect 476204 708678 476804 709670
rect 476204 708442 476386 708678
rect 476622 708442 476804 708678
rect 476204 708358 476804 708442
rect 476204 708122 476386 708358
rect 476622 708122 476804 708358
rect 472504 706758 473104 707750
rect 472504 706522 472686 706758
rect 472922 706522 473104 706758
rect 472504 706438 473104 706522
rect 472504 706202 472686 706438
rect 472922 706202 473104 706438
rect 461904 679158 462086 679394
rect 462322 679158 462504 679394
rect 461904 643394 462504 679158
rect 461904 643158 462086 643394
rect 462322 643158 462504 643394
rect 461904 607394 462504 643158
rect 461904 607158 462086 607394
rect 462322 607158 462504 607394
rect 461904 571394 462504 607158
rect 461904 571158 462086 571394
rect 462322 571158 462504 571394
rect 461904 535394 462504 571158
rect 461904 535158 462086 535394
rect 462322 535158 462504 535394
rect 461904 499394 462504 535158
rect 461904 499158 462086 499394
rect 462322 499158 462504 499394
rect 461904 463394 462504 499158
rect 461904 463158 462086 463394
rect 462322 463158 462504 463394
rect 461904 427394 462504 463158
rect 461904 427158 462086 427394
rect 462322 427158 462504 427394
rect 461904 425308 462504 427158
rect 468804 704838 469404 705830
rect 468804 704602 468986 704838
rect 469222 704602 469404 704838
rect 468804 704518 469404 704602
rect 468804 704282 468986 704518
rect 469222 704282 469404 704518
rect 468804 686294 469404 704282
rect 468804 686058 468986 686294
rect 469222 686058 469404 686294
rect 468804 650294 469404 686058
rect 468804 650058 468986 650294
rect 469222 650058 469404 650294
rect 468804 614294 469404 650058
rect 468804 614058 468986 614294
rect 469222 614058 469404 614294
rect 468804 578294 469404 614058
rect 468804 578058 468986 578294
rect 469222 578058 469404 578294
rect 468804 542294 469404 578058
rect 468804 542058 468986 542294
rect 469222 542058 469404 542294
rect 468804 506294 469404 542058
rect 468804 506058 468986 506294
rect 469222 506058 469404 506294
rect 468804 470294 469404 506058
rect 468804 470058 468986 470294
rect 469222 470058 469404 470294
rect 468804 434294 469404 470058
rect 468804 434058 468986 434294
rect 469222 434058 469404 434294
rect 468804 425308 469404 434058
rect 472504 689994 473104 706202
rect 472504 689758 472686 689994
rect 472922 689758 473104 689994
rect 472504 653994 473104 689758
rect 472504 653758 472686 653994
rect 472922 653758 473104 653994
rect 472504 617994 473104 653758
rect 472504 617758 472686 617994
rect 472922 617758 473104 617994
rect 472504 581994 473104 617758
rect 472504 581758 472686 581994
rect 472922 581758 473104 581994
rect 472504 545994 473104 581758
rect 472504 545758 472686 545994
rect 472922 545758 473104 545994
rect 472504 509994 473104 545758
rect 472504 509758 472686 509994
rect 472922 509758 473104 509994
rect 472504 473994 473104 509758
rect 472504 473758 472686 473994
rect 472922 473758 473104 473994
rect 472504 437994 473104 473758
rect 472504 437758 472686 437994
rect 472922 437758 473104 437994
rect 472504 425308 473104 437758
rect 476204 693694 476804 708122
rect 476204 693458 476386 693694
rect 476622 693458 476804 693694
rect 476204 657694 476804 693458
rect 476204 657458 476386 657694
rect 476622 657458 476804 657694
rect 476204 621694 476804 657458
rect 476204 621458 476386 621694
rect 476622 621458 476804 621694
rect 476204 585694 476804 621458
rect 476204 585458 476386 585694
rect 476622 585458 476804 585694
rect 476204 549694 476804 585458
rect 476204 549458 476386 549694
rect 476622 549458 476804 549694
rect 476204 513694 476804 549458
rect 476204 513458 476386 513694
rect 476622 513458 476804 513694
rect 476204 477694 476804 513458
rect 476204 477458 476386 477694
rect 476622 477458 476804 477694
rect 476204 441694 476804 477458
rect 476204 441458 476386 441694
rect 476622 441458 476804 441694
rect 476204 425308 476804 441458
rect 479904 697394 480504 710042
rect 497904 711558 498504 711590
rect 497904 711322 498086 711558
rect 498322 711322 498504 711558
rect 497904 711238 498504 711322
rect 497904 711002 498086 711238
rect 498322 711002 498504 711238
rect 494204 709638 494804 709670
rect 494204 709402 494386 709638
rect 494622 709402 494804 709638
rect 494204 709318 494804 709402
rect 494204 709082 494386 709318
rect 494622 709082 494804 709318
rect 490504 707718 491104 707750
rect 490504 707482 490686 707718
rect 490922 707482 491104 707718
rect 490504 707398 491104 707482
rect 490504 707162 490686 707398
rect 490922 707162 491104 707398
rect 479904 697158 480086 697394
rect 480322 697158 480504 697394
rect 479904 661394 480504 697158
rect 479904 661158 480086 661394
rect 480322 661158 480504 661394
rect 479904 625394 480504 661158
rect 479904 625158 480086 625394
rect 480322 625158 480504 625394
rect 479904 589394 480504 625158
rect 479904 589158 480086 589394
rect 480322 589158 480504 589394
rect 479904 553394 480504 589158
rect 479904 553158 480086 553394
rect 480322 553158 480504 553394
rect 479904 517394 480504 553158
rect 479904 517158 480086 517394
rect 480322 517158 480504 517394
rect 479904 481394 480504 517158
rect 479904 481158 480086 481394
rect 480322 481158 480504 481394
rect 479904 445394 480504 481158
rect 479904 445158 480086 445394
rect 480322 445158 480504 445394
rect 340272 416294 340620 416476
rect 340272 416058 340328 416294
rect 340564 416058 340620 416294
rect 340272 415876 340620 416058
rect 476000 416294 476348 416476
rect 476000 416058 476056 416294
rect 476292 416058 476348 416294
rect 476000 415876 476348 416058
rect 335904 409158 336086 409394
rect 336322 409158 336504 409394
rect 335904 373394 336504 409158
rect 479904 409394 480504 445158
rect 479904 409158 480086 409394
rect 480322 409158 480504 409394
rect 340952 398294 341300 398476
rect 340952 398058 341008 398294
rect 341244 398058 341300 398294
rect 340952 397876 341300 398058
rect 475320 398294 475668 398476
rect 475320 398058 475376 398294
rect 475612 398058 475668 398294
rect 475320 397876 475668 398058
rect 340272 380294 340620 380476
rect 340272 380058 340328 380294
rect 340564 380058 340620 380294
rect 340272 379876 340620 380058
rect 476000 380294 476348 380476
rect 476000 380058 476056 380294
rect 476292 380058 476348 380294
rect 476000 379876 476348 380058
rect 335904 373158 336086 373394
rect 336322 373158 336504 373394
rect 335904 337394 336504 373158
rect 479904 373394 480504 409158
rect 479904 373158 480086 373394
rect 480322 373158 480504 373394
rect 340952 362294 341300 362476
rect 340952 362058 341008 362294
rect 341244 362058 341300 362294
rect 340952 361876 341300 362058
rect 475320 362294 475668 362476
rect 475320 362058 475376 362294
rect 475612 362058 475668 362294
rect 475320 361876 475668 362058
rect 340272 344294 340620 344476
rect 340272 344058 340328 344294
rect 340564 344058 340620 344294
rect 340272 343876 340620 344058
rect 476000 344294 476348 344476
rect 476000 344058 476056 344294
rect 476292 344058 476348 344294
rect 476000 343876 476348 344058
rect 393454 340076 393622 340136
rect 356056 339690 356116 340000
rect 357144 339690 357204 340000
rect 358232 339690 358292 340000
rect 356056 339630 356162 339690
rect 335904 337158 336086 337394
rect 336322 337158 336504 337394
rect 335904 301394 336504 337158
rect 335904 301158 336086 301394
rect 336322 301158 336504 301394
rect 335904 265394 336504 301158
rect 335904 265158 336086 265394
rect 336322 265158 336504 265394
rect 335904 229394 336504 265158
rect 335904 229158 336086 229394
rect 336322 229158 336504 229394
rect 335904 193394 336504 229158
rect 335904 193158 336086 193394
rect 336322 193158 336504 193394
rect 335904 157394 336504 193158
rect 335904 157158 336086 157394
rect 336322 157158 336504 157394
rect 335904 121394 336504 157158
rect 335904 121158 336086 121394
rect 336322 121158 336504 121394
rect 335904 85394 336504 121158
rect 335904 85158 336086 85394
rect 336322 85158 336504 85394
rect 335904 49394 336504 85158
rect 335904 49158 336086 49394
rect 336322 49158 336504 49394
rect 335904 13394 336504 49158
rect 335904 13158 336086 13394
rect 336322 13158 336504 13394
rect 317904 -7302 318086 -7066
rect 318322 -7302 318504 -7066
rect 317904 -7386 318504 -7302
rect 317904 -7622 318086 -7386
rect 318322 -7622 318504 -7386
rect 317904 -7654 318504 -7622
rect 335904 -6106 336504 13158
rect 342804 308294 343404 338000
rect 342804 308058 342986 308294
rect 343222 308058 343404 308294
rect 342804 272294 343404 308058
rect 342804 272058 342986 272294
rect 343222 272058 343404 272294
rect 342804 236294 343404 272058
rect 342804 236058 342986 236294
rect 343222 236058 343404 236294
rect 342804 200294 343404 236058
rect 342804 200058 342986 200294
rect 343222 200058 343404 200294
rect 342804 164294 343404 200058
rect 342804 164058 342986 164294
rect 343222 164058 343404 164294
rect 342804 128294 343404 164058
rect 342804 128058 342986 128294
rect 343222 128058 343404 128294
rect 342804 92294 343404 128058
rect 342804 92058 342986 92294
rect 343222 92058 343404 92294
rect 342804 56294 343404 92058
rect 342804 56058 342986 56294
rect 343222 56058 343404 56294
rect 342804 20294 343404 56058
rect 342804 20058 342986 20294
rect 343222 20058 343404 20294
rect 342804 -1306 343404 20058
rect 342804 -1542 342986 -1306
rect 343222 -1542 343404 -1306
rect 342804 -1626 343404 -1542
rect 342804 -1862 342986 -1626
rect 343222 -1862 343404 -1626
rect 342804 -1894 343404 -1862
rect 346504 311994 347104 338000
rect 346504 311758 346686 311994
rect 346922 311758 347104 311994
rect 346504 275994 347104 311758
rect 346504 275758 346686 275994
rect 346922 275758 347104 275994
rect 346504 239994 347104 275758
rect 346504 239758 346686 239994
rect 346922 239758 347104 239994
rect 346504 203994 347104 239758
rect 346504 203758 346686 203994
rect 346922 203758 347104 203994
rect 346504 167994 347104 203758
rect 346504 167758 346686 167994
rect 346922 167758 347104 167994
rect 346504 131994 347104 167758
rect 346504 131758 346686 131994
rect 346922 131758 347104 131994
rect 346504 95994 347104 131758
rect 346504 95758 346686 95994
rect 346922 95758 347104 95994
rect 346504 59994 347104 95758
rect 346504 59758 346686 59994
rect 346922 59758 347104 59994
rect 346504 23994 347104 59758
rect 346504 23758 346686 23994
rect 346922 23758 347104 23994
rect 346504 -3226 347104 23758
rect 346504 -3462 346686 -3226
rect 346922 -3462 347104 -3226
rect 346504 -3546 347104 -3462
rect 346504 -3782 346686 -3546
rect 346922 -3782 347104 -3546
rect 346504 -3814 347104 -3782
rect 350204 315694 350804 338000
rect 350204 315458 350386 315694
rect 350622 315458 350804 315694
rect 350204 279694 350804 315458
rect 350204 279458 350386 279694
rect 350622 279458 350804 279694
rect 350204 243694 350804 279458
rect 350204 243458 350386 243694
rect 350622 243458 350804 243694
rect 350204 207694 350804 243458
rect 350204 207458 350386 207694
rect 350622 207458 350804 207694
rect 350204 171694 350804 207458
rect 350204 171458 350386 171694
rect 350622 171458 350804 171694
rect 350204 135694 350804 171458
rect 350204 135458 350386 135694
rect 350622 135458 350804 135694
rect 350204 99694 350804 135458
rect 350204 99458 350386 99694
rect 350622 99458 350804 99694
rect 350204 63694 350804 99458
rect 350204 63458 350386 63694
rect 350622 63458 350804 63694
rect 350204 27694 350804 63458
rect 350204 27458 350386 27694
rect 350622 27458 350804 27694
rect 350204 -5146 350804 27458
rect 350204 -5382 350386 -5146
rect 350622 -5382 350804 -5146
rect 350204 -5466 350804 -5382
rect 350204 -5702 350386 -5466
rect 350622 -5702 350804 -5466
rect 350204 -5734 350804 -5702
rect 353904 319394 354504 338000
rect 356102 337381 356162 339630
rect 357022 339630 357204 339690
rect 358126 339630 358292 339690
rect 359592 339690 359652 340000
rect 360544 339690 360604 340000
rect 359592 339630 359658 339690
rect 357022 337653 357082 339630
rect 358126 337653 358186 339630
rect 359598 337653 359658 339630
rect 360518 339630 360604 339690
rect 361768 339690 361828 340000
rect 363128 339690 363188 340000
rect 364216 339690 364276 340000
rect 361768 339630 361866 339690
rect 360518 337653 360578 339630
rect 357019 337652 357085 337653
rect 357019 337588 357020 337652
rect 357084 337588 357085 337652
rect 357019 337587 357085 337588
rect 358123 337652 358189 337653
rect 358123 337588 358124 337652
rect 358188 337588 358189 337652
rect 358123 337587 358189 337588
rect 359595 337652 359661 337653
rect 359595 337588 359596 337652
rect 359660 337588 359661 337652
rect 359595 337587 359661 337588
rect 360515 337652 360581 337653
rect 360515 337588 360516 337652
rect 360580 337588 360581 337652
rect 360515 337587 360581 337588
rect 356099 337380 356165 337381
rect 356099 337316 356100 337380
rect 356164 337316 356165 337380
rect 356099 337315 356165 337316
rect 353904 319158 354086 319394
rect 354322 319158 354504 319394
rect 353904 283394 354504 319158
rect 353904 283158 354086 283394
rect 354322 283158 354504 283394
rect 353904 247394 354504 283158
rect 353904 247158 354086 247394
rect 354322 247158 354504 247394
rect 353904 211394 354504 247158
rect 353904 211158 354086 211394
rect 354322 211158 354504 211394
rect 353904 175394 354504 211158
rect 353904 175158 354086 175394
rect 354322 175158 354504 175394
rect 353904 139394 354504 175158
rect 353904 139158 354086 139394
rect 354322 139158 354504 139394
rect 353904 103394 354504 139158
rect 353904 103158 354086 103394
rect 354322 103158 354504 103394
rect 353904 67394 354504 103158
rect 353904 67158 354086 67394
rect 354322 67158 354504 67394
rect 353904 31394 354504 67158
rect 353904 31158 354086 31394
rect 354322 31158 354504 31394
rect 335904 -6342 336086 -6106
rect 336322 -6342 336504 -6106
rect 335904 -6426 336504 -6342
rect 335904 -6662 336086 -6426
rect 336322 -6662 336504 -6426
rect 335904 -7654 336504 -6662
rect 353904 -7066 354504 31158
rect 360804 326294 361404 338000
rect 361806 337653 361866 339630
rect 363094 339630 363188 339690
rect 364198 339630 364276 339690
rect 363094 337653 363154 339630
rect 364198 337789 364258 339630
rect 365440 339510 365500 340000
rect 366528 339510 366588 340000
rect 367616 339510 367676 340000
rect 368296 339510 368356 340000
rect 365440 339450 365546 339510
rect 364195 337788 364261 337789
rect 364195 337724 364196 337788
rect 364260 337724 364261 337788
rect 364195 337723 364261 337724
rect 361803 337652 361869 337653
rect 361803 337588 361804 337652
rect 361868 337588 361869 337652
rect 361803 337587 361869 337588
rect 363091 337652 363157 337653
rect 363091 337588 363092 337652
rect 363156 337588 363157 337652
rect 363091 337587 363157 337588
rect 360804 326058 360986 326294
rect 361222 326058 361404 326294
rect 360804 290294 361404 326058
rect 360804 290058 360986 290294
rect 361222 290058 361404 290294
rect 360804 254294 361404 290058
rect 360804 254058 360986 254294
rect 361222 254058 361404 254294
rect 360804 218294 361404 254058
rect 360804 218058 360986 218294
rect 361222 218058 361404 218294
rect 360804 182294 361404 218058
rect 360804 182058 360986 182294
rect 361222 182058 361404 182294
rect 360804 146294 361404 182058
rect 360804 146058 360986 146294
rect 361222 146058 361404 146294
rect 360804 110294 361404 146058
rect 360804 110058 360986 110294
rect 361222 110058 361404 110294
rect 360804 74294 361404 110058
rect 360804 74058 360986 74294
rect 361222 74058 361404 74294
rect 360804 38294 361404 74058
rect 360804 38058 360986 38294
rect 361222 38058 361404 38294
rect 360804 2294 361404 38058
rect 360804 2058 360986 2294
rect 361222 2058 361404 2294
rect 360804 -346 361404 2058
rect 360804 -582 360986 -346
rect 361222 -582 361404 -346
rect 360804 -666 361404 -582
rect 360804 -902 360986 -666
rect 361222 -902 361404 -666
rect 360804 -1894 361404 -902
rect 364504 329994 365104 338000
rect 365486 336837 365546 339450
rect 366406 339450 366588 339510
rect 367510 339450 367676 339510
rect 368062 339450 368356 339510
rect 368704 339510 368764 340000
rect 370064 339510 370124 340000
rect 370744 339510 370804 340000
rect 371288 339510 371348 340000
rect 372376 339510 372436 340000
rect 373464 339690 373524 340000
rect 368704 339450 369042 339510
rect 370064 339450 370146 339510
rect 366406 337653 366466 339450
rect 367510 337789 367570 339450
rect 367507 337788 367573 337789
rect 367507 337724 367508 337788
rect 367572 337724 367573 337788
rect 367507 337723 367573 337724
rect 368062 337653 368122 339450
rect 366403 337652 366469 337653
rect 366403 337588 366404 337652
rect 366468 337588 366469 337652
rect 366403 337587 366469 337588
rect 368059 337652 368125 337653
rect 368059 337588 368060 337652
rect 368124 337588 368125 337652
rect 368059 337587 368125 337588
rect 365483 336836 365549 336837
rect 365483 336772 365484 336836
rect 365548 336772 365549 336836
rect 365483 336771 365549 336772
rect 364504 329758 364686 329994
rect 364922 329758 365104 329994
rect 364504 293994 365104 329758
rect 364504 293758 364686 293994
rect 364922 293758 365104 293994
rect 364504 257994 365104 293758
rect 364504 257758 364686 257994
rect 364922 257758 365104 257994
rect 364504 221994 365104 257758
rect 364504 221758 364686 221994
rect 364922 221758 365104 221994
rect 364504 185994 365104 221758
rect 364504 185758 364686 185994
rect 364922 185758 365104 185994
rect 364504 149994 365104 185758
rect 364504 149758 364686 149994
rect 364922 149758 365104 149994
rect 364504 113994 365104 149758
rect 364504 113758 364686 113994
rect 364922 113758 365104 113994
rect 364504 77994 365104 113758
rect 364504 77758 364686 77994
rect 364922 77758 365104 77994
rect 364504 41994 365104 77758
rect 364504 41758 364686 41994
rect 364922 41758 365104 41994
rect 364504 5994 365104 41758
rect 364504 5758 364686 5994
rect 364922 5758 365104 5994
rect 364504 -2266 365104 5758
rect 364504 -2502 364686 -2266
rect 364922 -2502 365104 -2266
rect 364504 -2586 365104 -2502
rect 364504 -2822 364686 -2586
rect 364922 -2822 365104 -2586
rect 364504 -3814 365104 -2822
rect 368204 333694 368804 338000
rect 368982 337653 369042 339450
rect 370086 337789 370146 339450
rect 370638 339450 370804 339510
rect 371190 339450 371348 339510
rect 372294 339450 372436 339510
rect 373398 339630 373524 339690
rect 370083 337788 370149 337789
rect 370083 337724 370084 337788
rect 370148 337724 370149 337788
rect 370083 337723 370149 337724
rect 370638 337653 370698 339450
rect 368979 337652 369045 337653
rect 368979 337588 368980 337652
rect 369044 337588 369045 337652
rect 368979 337587 369045 337588
rect 370635 337652 370701 337653
rect 370635 337588 370636 337652
rect 370700 337588 370701 337652
rect 370635 337587 370701 337588
rect 371190 336837 371250 339450
rect 372294 338197 372354 339450
rect 372291 338196 372357 338197
rect 372291 338132 372292 338196
rect 372356 338132 372357 338196
rect 372291 338131 372357 338132
rect 371904 337394 372504 338000
rect 373398 337653 373458 339630
rect 373600 339510 373660 340000
rect 374552 339510 374612 340000
rect 375912 339510 375972 340000
rect 373582 339450 373660 339510
rect 374502 339450 374612 339510
rect 375790 339450 375972 339510
rect 376048 339510 376108 340000
rect 377000 339510 377060 340000
rect 378088 339510 378148 340000
rect 376048 339450 376218 339510
rect 373582 337789 373642 339450
rect 373579 337788 373645 337789
rect 373579 337724 373580 337788
rect 373644 337724 373645 337788
rect 373579 337723 373645 337724
rect 374502 337653 374562 339450
rect 375790 337653 375850 339450
rect 376158 337925 376218 339450
rect 376894 339450 377060 339510
rect 377998 339450 378148 339510
rect 378496 339510 378556 340000
rect 379448 339690 379508 340000
rect 379448 339630 379530 339690
rect 378496 339450 378610 339510
rect 376155 337924 376221 337925
rect 376155 337860 376156 337924
rect 376220 337860 376221 337924
rect 376155 337859 376221 337860
rect 373395 337652 373461 337653
rect 373395 337588 373396 337652
rect 373460 337588 373461 337652
rect 373395 337587 373461 337588
rect 374499 337652 374565 337653
rect 374499 337588 374500 337652
rect 374564 337588 374565 337652
rect 374499 337587 374565 337588
rect 375787 337652 375853 337653
rect 375787 337588 375788 337652
rect 375852 337588 375853 337652
rect 375787 337587 375853 337588
rect 371904 337158 372086 337394
rect 372322 337158 372504 337394
rect 371187 336836 371253 336837
rect 371187 336772 371188 336836
rect 371252 336772 371253 336836
rect 371187 336771 371253 336772
rect 368204 333458 368386 333694
rect 368622 333458 368804 333694
rect 368204 297694 368804 333458
rect 368204 297458 368386 297694
rect 368622 297458 368804 297694
rect 368204 261694 368804 297458
rect 368204 261458 368386 261694
rect 368622 261458 368804 261694
rect 368204 225694 368804 261458
rect 368204 225458 368386 225694
rect 368622 225458 368804 225694
rect 368204 189694 368804 225458
rect 368204 189458 368386 189694
rect 368622 189458 368804 189694
rect 368204 153694 368804 189458
rect 368204 153458 368386 153694
rect 368622 153458 368804 153694
rect 368204 117694 368804 153458
rect 368204 117458 368386 117694
rect 368622 117458 368804 117694
rect 368204 81694 368804 117458
rect 368204 81458 368386 81694
rect 368622 81458 368804 81694
rect 368204 45694 368804 81458
rect 368204 45458 368386 45694
rect 368622 45458 368804 45694
rect 368204 9694 368804 45458
rect 368204 9458 368386 9694
rect 368622 9458 368804 9694
rect 368204 -4186 368804 9458
rect 368204 -4422 368386 -4186
rect 368622 -4422 368804 -4186
rect 368204 -4506 368804 -4422
rect 368204 -4742 368386 -4506
rect 368622 -4742 368804 -4506
rect 368204 -5734 368804 -4742
rect 371904 301394 372504 337158
rect 376894 336837 376954 339450
rect 377998 337653 378058 339450
rect 378550 337789 378610 339450
rect 378547 337788 378613 337789
rect 378547 337724 378548 337788
rect 378612 337724 378613 337788
rect 378547 337723 378613 337724
rect 377995 337652 378061 337653
rect 377995 337588 377996 337652
rect 378060 337588 378061 337652
rect 377995 337587 378061 337588
rect 376891 336836 376957 336837
rect 376891 336772 376892 336836
rect 376956 336772 376957 336836
rect 376891 336771 376957 336772
rect 371904 301158 372086 301394
rect 372322 301158 372504 301394
rect 371904 265394 372504 301158
rect 371904 265158 372086 265394
rect 372322 265158 372504 265394
rect 371904 229394 372504 265158
rect 371904 229158 372086 229394
rect 372322 229158 372504 229394
rect 371904 193394 372504 229158
rect 371904 193158 372086 193394
rect 372322 193158 372504 193394
rect 371904 157394 372504 193158
rect 371904 157158 372086 157394
rect 372322 157158 372504 157394
rect 371904 121394 372504 157158
rect 371904 121158 372086 121394
rect 372322 121158 372504 121394
rect 371904 85394 372504 121158
rect 371904 85158 372086 85394
rect 372322 85158 372504 85394
rect 371904 49394 372504 85158
rect 371904 49158 372086 49394
rect 372322 49158 372504 49394
rect 371904 13394 372504 49158
rect 371904 13158 372086 13394
rect 372322 13158 372504 13394
rect 353904 -7302 354086 -7066
rect 354322 -7302 354504 -7066
rect 353904 -7386 354504 -7302
rect 353904 -7622 354086 -7386
rect 354322 -7622 354504 -7386
rect 353904 -7654 354504 -7622
rect 371904 -6106 372504 13158
rect 378804 308294 379404 338000
rect 379470 337925 379530 339630
rect 380672 339510 380732 340000
rect 380574 339450 380732 339510
rect 381080 339510 381140 340000
rect 381760 339510 381820 340000
rect 382848 339510 382908 340000
rect 383528 339510 383588 340000
rect 383936 339510 383996 340000
rect 385296 339510 385356 340000
rect 385976 339510 386036 340000
rect 381080 339450 381186 339510
rect 379467 337924 379533 337925
rect 379467 337860 379468 337924
rect 379532 337860 379533 337924
rect 379467 337859 379533 337860
rect 380574 337109 380634 339450
rect 381126 337653 381186 339450
rect 381678 339450 381820 339510
rect 382782 339450 382908 339510
rect 383518 339450 383588 339510
rect 383886 339450 383996 339510
rect 385174 339450 385356 339510
rect 385910 339450 386036 339510
rect 386384 339510 386444 340000
rect 387608 339510 387668 340000
rect 386384 339450 386522 339510
rect 381678 337789 381738 339450
rect 382782 338197 382842 339450
rect 382779 338196 382845 338197
rect 382779 338132 382780 338196
rect 382844 338132 382845 338196
rect 382779 338131 382845 338132
rect 381675 337788 381741 337789
rect 381675 337724 381676 337788
rect 381740 337724 381741 337788
rect 381675 337723 381741 337724
rect 381123 337652 381189 337653
rect 381123 337588 381124 337652
rect 381188 337588 381189 337652
rect 381123 337587 381189 337588
rect 380571 337108 380637 337109
rect 380571 337044 380572 337108
rect 380636 337044 380637 337108
rect 380571 337043 380637 337044
rect 378804 308058 378986 308294
rect 379222 308058 379404 308294
rect 378804 272294 379404 308058
rect 378804 272058 378986 272294
rect 379222 272058 379404 272294
rect 378804 236294 379404 272058
rect 378804 236058 378986 236294
rect 379222 236058 379404 236294
rect 378804 200294 379404 236058
rect 378804 200058 378986 200294
rect 379222 200058 379404 200294
rect 378804 164294 379404 200058
rect 378804 164058 378986 164294
rect 379222 164058 379404 164294
rect 378804 128294 379404 164058
rect 378804 128058 378986 128294
rect 379222 128058 379404 128294
rect 378804 92294 379404 128058
rect 378804 92058 378986 92294
rect 379222 92058 379404 92294
rect 378804 56294 379404 92058
rect 378804 56058 378986 56294
rect 379222 56058 379404 56294
rect 378804 20294 379404 56058
rect 378804 20058 378986 20294
rect 379222 20058 379404 20294
rect 378804 -1306 379404 20058
rect 378804 -1542 378986 -1306
rect 379222 -1542 379404 -1306
rect 378804 -1626 379404 -1542
rect 378804 -1862 378986 -1626
rect 379222 -1862 379404 -1626
rect 378804 -1894 379404 -1862
rect 382504 311994 383104 338000
rect 383518 337381 383578 339450
rect 383515 337380 383581 337381
rect 383515 337316 383516 337380
rect 383580 337316 383581 337380
rect 383515 337315 383581 337316
rect 383886 336973 383946 339450
rect 385174 337653 385234 339450
rect 385171 337652 385237 337653
rect 385171 337588 385172 337652
rect 385236 337588 385237 337652
rect 385171 337587 385237 337588
rect 385910 337517 385970 339450
rect 386462 338197 386522 339450
rect 387566 339450 387668 339510
rect 388288 339510 388348 340000
rect 388696 339510 388756 340000
rect 389784 339510 389844 340000
rect 388288 339450 388362 339510
rect 386459 338196 386525 338197
rect 386459 338132 386460 338196
rect 386524 338132 386525 338196
rect 386459 338131 386525 338132
rect 385907 337516 385973 337517
rect 385907 337452 385908 337516
rect 385972 337452 385973 337516
rect 385907 337451 385973 337452
rect 383883 336972 383949 336973
rect 383883 336908 383884 336972
rect 383948 336908 383949 336972
rect 383883 336907 383949 336908
rect 382504 311758 382686 311994
rect 382922 311758 383104 311994
rect 382504 275994 383104 311758
rect 382504 275758 382686 275994
rect 382922 275758 383104 275994
rect 382504 239994 383104 275758
rect 382504 239758 382686 239994
rect 382922 239758 383104 239994
rect 382504 203994 383104 239758
rect 382504 203758 382686 203994
rect 382922 203758 383104 203994
rect 382504 167994 383104 203758
rect 382504 167758 382686 167994
rect 382922 167758 383104 167994
rect 382504 131994 383104 167758
rect 382504 131758 382686 131994
rect 382922 131758 383104 131994
rect 382504 95994 383104 131758
rect 382504 95758 382686 95994
rect 382922 95758 383104 95994
rect 382504 59994 383104 95758
rect 382504 59758 382686 59994
rect 382922 59758 383104 59994
rect 382504 23994 383104 59758
rect 382504 23758 382686 23994
rect 382922 23758 383104 23994
rect 382504 -3226 383104 23758
rect 382504 -3462 382686 -3226
rect 382922 -3462 383104 -3226
rect 382504 -3546 383104 -3462
rect 382504 -3782 382686 -3546
rect 382922 -3782 383104 -3546
rect 382504 -3814 383104 -3782
rect 386204 315694 386804 338000
rect 387566 337245 387626 339450
rect 388302 337517 388362 339450
rect 388670 339450 388756 339510
rect 389774 339450 389844 339510
rect 391008 339510 391068 340000
rect 391144 339690 391204 340000
rect 391144 339630 391306 339690
rect 391008 339450 391122 339510
rect 388299 337516 388365 337517
rect 388299 337452 388300 337516
rect 388364 337452 388365 337516
rect 388299 337451 388365 337452
rect 387563 337244 387629 337245
rect 387563 337180 387564 337244
rect 387628 337180 387629 337244
rect 387563 337179 387629 337180
rect 388670 337109 388730 339450
rect 389774 337789 389834 339450
rect 389771 337788 389837 337789
rect 389771 337724 389772 337788
rect 389836 337724 389837 337788
rect 389771 337723 389837 337724
rect 388667 337108 388733 337109
rect 388667 337044 388668 337108
rect 388732 337044 388733 337108
rect 388667 337043 388733 337044
rect 386204 315458 386386 315694
rect 386622 315458 386804 315694
rect 386204 279694 386804 315458
rect 386204 279458 386386 279694
rect 386622 279458 386804 279694
rect 386204 243694 386804 279458
rect 386204 243458 386386 243694
rect 386622 243458 386804 243694
rect 386204 207694 386804 243458
rect 386204 207458 386386 207694
rect 386622 207458 386804 207694
rect 386204 171694 386804 207458
rect 386204 171458 386386 171694
rect 386622 171458 386804 171694
rect 386204 135694 386804 171458
rect 386204 135458 386386 135694
rect 386622 135458 386804 135694
rect 386204 99694 386804 135458
rect 386204 99458 386386 99694
rect 386622 99458 386804 99694
rect 386204 63694 386804 99458
rect 386204 63458 386386 63694
rect 386622 63458 386804 63694
rect 386204 27694 386804 63458
rect 386204 27458 386386 27694
rect 386622 27458 386804 27694
rect 386204 -5146 386804 27458
rect 386204 -5382 386386 -5146
rect 386622 -5382 386804 -5146
rect 386204 -5466 386804 -5382
rect 386204 -5702 386386 -5466
rect 386622 -5702 386804 -5466
rect 386204 -5734 386804 -5702
rect 389904 319394 390504 338000
rect 391062 337653 391122 339450
rect 391059 337652 391125 337653
rect 391059 337588 391060 337652
rect 391124 337588 391125 337652
rect 391059 337587 391125 337588
rect 391246 336837 391306 339630
rect 392232 339510 392292 340000
rect 393320 339690 393380 340000
rect 392166 339450 392292 339510
rect 393086 339630 393380 339690
rect 392166 337789 392226 339450
rect 392163 337788 392229 337789
rect 392163 337724 392164 337788
rect 392228 337724 392229 337788
rect 392163 337723 392229 337724
rect 393086 336973 393146 339630
rect 393454 337653 393514 340076
rect 394408 339690 394468 340000
rect 395768 339690 395828 340000
rect 396040 339690 396100 340000
rect 396992 339690 397052 340000
rect 398080 339690 398140 340000
rect 398488 339690 398548 340000
rect 399168 339690 399228 340000
rect 394374 339630 394468 339690
rect 395662 339630 395828 339690
rect 396030 339630 396100 339690
rect 396582 339630 397052 339690
rect 398054 339630 398140 339690
rect 398422 339630 398548 339690
rect 399158 339630 399228 339690
rect 400936 339690 400996 340000
rect 403520 339690 403580 340000
rect 405968 339690 406028 340000
rect 408280 339690 408340 340000
rect 411000 339690 411060 340000
rect 413448 339690 413508 340000
rect 400936 339630 401242 339690
rect 403520 339630 403634 339690
rect 393451 337652 393517 337653
rect 393451 337588 393452 337652
rect 393516 337588 393517 337652
rect 393451 337587 393517 337588
rect 394374 337109 394434 339630
rect 395662 337925 395722 339630
rect 395659 337924 395725 337925
rect 395659 337860 395660 337924
rect 395724 337860 395725 337924
rect 395659 337859 395725 337860
rect 396030 337653 396090 339630
rect 396027 337652 396093 337653
rect 396027 337588 396028 337652
rect 396092 337588 396093 337652
rect 396027 337587 396093 337588
rect 394371 337108 394437 337109
rect 394371 337044 394372 337108
rect 394436 337044 394437 337108
rect 394371 337043 394437 337044
rect 396582 336973 396642 339630
rect 393083 336972 393149 336973
rect 393083 336908 393084 336972
rect 393148 336908 393149 336972
rect 393083 336907 393149 336908
rect 396579 336972 396645 336973
rect 396579 336908 396580 336972
rect 396644 336908 396645 336972
rect 396579 336907 396645 336908
rect 391243 336836 391309 336837
rect 391243 336772 391244 336836
rect 391308 336772 391309 336836
rect 391243 336771 391309 336772
rect 389904 319158 390086 319394
rect 390322 319158 390504 319394
rect 389904 283394 390504 319158
rect 389904 283158 390086 283394
rect 390322 283158 390504 283394
rect 389904 247394 390504 283158
rect 389904 247158 390086 247394
rect 390322 247158 390504 247394
rect 389904 211394 390504 247158
rect 389904 211158 390086 211394
rect 390322 211158 390504 211394
rect 389904 175394 390504 211158
rect 389904 175158 390086 175394
rect 390322 175158 390504 175394
rect 389904 139394 390504 175158
rect 389904 139158 390086 139394
rect 390322 139158 390504 139394
rect 389904 103394 390504 139158
rect 389904 103158 390086 103394
rect 390322 103158 390504 103394
rect 389904 67394 390504 103158
rect 389904 67158 390086 67394
rect 390322 67158 390504 67394
rect 389904 31394 390504 67158
rect 389904 31158 390086 31394
rect 390322 31158 390504 31394
rect 371904 -6342 372086 -6106
rect 372322 -6342 372504 -6106
rect 371904 -6426 372504 -6342
rect 371904 -6662 372086 -6426
rect 372322 -6662 372504 -6426
rect 371904 -7654 372504 -6662
rect 389904 -7066 390504 31158
rect 396804 326294 397404 338000
rect 398054 337925 398114 339630
rect 398051 337924 398117 337925
rect 398051 337860 398052 337924
rect 398116 337860 398117 337924
rect 398051 337859 398117 337860
rect 398422 336837 398482 339630
rect 399158 337653 399218 339630
rect 399155 337652 399221 337653
rect 399155 337588 399156 337652
rect 399220 337588 399221 337652
rect 399155 337587 399221 337588
rect 398419 336836 398485 336837
rect 398419 336772 398420 336836
rect 398484 336772 398485 336836
rect 398419 336771 398485 336772
rect 396804 326058 396986 326294
rect 397222 326058 397404 326294
rect 396804 290294 397404 326058
rect 396804 290058 396986 290294
rect 397222 290058 397404 290294
rect 396804 254294 397404 290058
rect 396804 254058 396986 254294
rect 397222 254058 397404 254294
rect 396804 218294 397404 254058
rect 396804 218058 396986 218294
rect 397222 218058 397404 218294
rect 396804 182294 397404 218058
rect 396804 182058 396986 182294
rect 397222 182058 397404 182294
rect 396804 146294 397404 182058
rect 396804 146058 396986 146294
rect 397222 146058 397404 146294
rect 396804 110294 397404 146058
rect 396804 110058 396986 110294
rect 397222 110058 397404 110294
rect 396804 74294 397404 110058
rect 396804 74058 396986 74294
rect 397222 74058 397404 74294
rect 396804 38294 397404 74058
rect 396804 38058 396986 38294
rect 397222 38058 397404 38294
rect 396804 2294 397404 38058
rect 396804 2058 396986 2294
rect 397222 2058 397404 2294
rect 396804 -346 397404 2058
rect 396804 -582 396986 -346
rect 397222 -582 397404 -346
rect 396804 -666 397404 -582
rect 396804 -902 396986 -666
rect 397222 -902 397404 -666
rect 396804 -1894 397404 -902
rect 400504 329994 401104 338000
rect 401182 337653 401242 339630
rect 401179 337652 401245 337653
rect 401179 337588 401180 337652
rect 401244 337588 401245 337652
rect 401179 337587 401245 337588
rect 403574 336837 403634 339630
rect 405966 339630 406028 339690
rect 408174 339630 408340 339690
rect 410934 339630 411060 339690
rect 413326 339630 413508 339690
rect 415896 339690 415956 340000
rect 418480 339690 418540 340000
rect 420928 339690 420988 340000
rect 423512 339690 423572 340000
rect 425960 339690 426020 340000
rect 415896 339630 415962 339690
rect 403571 336836 403637 336837
rect 403571 336772 403572 336836
rect 403636 336772 403637 336836
rect 403571 336771 403637 336772
rect 400504 329758 400686 329994
rect 400922 329758 401104 329994
rect 400504 293994 401104 329758
rect 400504 293758 400686 293994
rect 400922 293758 401104 293994
rect 400504 257994 401104 293758
rect 400504 257758 400686 257994
rect 400922 257758 401104 257994
rect 400504 221994 401104 257758
rect 400504 221758 400686 221994
rect 400922 221758 401104 221994
rect 400504 185994 401104 221758
rect 400504 185758 400686 185994
rect 400922 185758 401104 185994
rect 400504 149994 401104 185758
rect 400504 149758 400686 149994
rect 400922 149758 401104 149994
rect 400504 113994 401104 149758
rect 400504 113758 400686 113994
rect 400922 113758 401104 113994
rect 400504 77994 401104 113758
rect 400504 77758 400686 77994
rect 400922 77758 401104 77994
rect 400504 41994 401104 77758
rect 400504 41758 400686 41994
rect 400922 41758 401104 41994
rect 400504 5994 401104 41758
rect 400504 5758 400686 5994
rect 400922 5758 401104 5994
rect 400504 -2266 401104 5758
rect 400504 -2502 400686 -2266
rect 400922 -2502 401104 -2266
rect 400504 -2586 401104 -2502
rect 400504 -2822 400686 -2586
rect 400922 -2822 401104 -2586
rect 400504 -3814 401104 -2822
rect 404204 333694 404804 338000
rect 405966 336973 406026 339630
rect 408174 338197 408234 339630
rect 408171 338196 408237 338197
rect 408171 338132 408172 338196
rect 408236 338132 408237 338196
rect 408171 338131 408237 338132
rect 407904 337394 408504 338000
rect 407904 337158 408086 337394
rect 408322 337158 408504 337394
rect 410934 337245 410994 339630
rect 413326 337653 413386 339630
rect 413323 337652 413389 337653
rect 413323 337588 413324 337652
rect 413388 337588 413389 337652
rect 413323 337587 413389 337588
rect 410931 337244 410997 337245
rect 410931 337180 410932 337244
rect 410996 337180 410997 337244
rect 410931 337179 410997 337180
rect 405963 336972 406029 336973
rect 405963 336908 405964 336972
rect 406028 336908 406029 336972
rect 405963 336907 406029 336908
rect 404204 333458 404386 333694
rect 404622 333458 404804 333694
rect 404204 297694 404804 333458
rect 404204 297458 404386 297694
rect 404622 297458 404804 297694
rect 404204 261694 404804 297458
rect 404204 261458 404386 261694
rect 404622 261458 404804 261694
rect 404204 225694 404804 261458
rect 404204 225458 404386 225694
rect 404622 225458 404804 225694
rect 404204 189694 404804 225458
rect 404204 189458 404386 189694
rect 404622 189458 404804 189694
rect 404204 153694 404804 189458
rect 404204 153458 404386 153694
rect 404622 153458 404804 153694
rect 404204 117694 404804 153458
rect 404204 117458 404386 117694
rect 404622 117458 404804 117694
rect 404204 81694 404804 117458
rect 404204 81458 404386 81694
rect 404622 81458 404804 81694
rect 404204 45694 404804 81458
rect 404204 45458 404386 45694
rect 404622 45458 404804 45694
rect 404204 9694 404804 45458
rect 404204 9458 404386 9694
rect 404622 9458 404804 9694
rect 404204 -4186 404804 9458
rect 404204 -4422 404386 -4186
rect 404622 -4422 404804 -4186
rect 404204 -4506 404804 -4422
rect 404204 -4742 404386 -4506
rect 404622 -4742 404804 -4506
rect 404204 -5734 404804 -4742
rect 407904 301394 408504 337158
rect 407904 301158 408086 301394
rect 408322 301158 408504 301394
rect 407904 265394 408504 301158
rect 407904 265158 408086 265394
rect 408322 265158 408504 265394
rect 407904 229394 408504 265158
rect 407904 229158 408086 229394
rect 408322 229158 408504 229394
rect 407904 193394 408504 229158
rect 407904 193158 408086 193394
rect 408322 193158 408504 193394
rect 407904 157394 408504 193158
rect 407904 157158 408086 157394
rect 408322 157158 408504 157394
rect 407904 121394 408504 157158
rect 407904 121158 408086 121394
rect 408322 121158 408504 121394
rect 407904 85394 408504 121158
rect 407904 85158 408086 85394
rect 408322 85158 408504 85394
rect 407904 49394 408504 85158
rect 407904 49158 408086 49394
rect 408322 49158 408504 49394
rect 407904 13394 408504 49158
rect 407904 13158 408086 13394
rect 408322 13158 408504 13394
rect 389904 -7302 390086 -7066
rect 390322 -7302 390504 -7066
rect 389904 -7386 390504 -7302
rect 389904 -7622 390086 -7386
rect 390322 -7622 390504 -7386
rect 389904 -7654 390504 -7622
rect 407904 -6106 408504 13158
rect 414804 308294 415404 338000
rect 415902 337653 415962 339630
rect 418294 339630 418540 339690
rect 420870 339630 420988 339690
rect 423446 339630 423572 339690
rect 425654 339630 426020 339690
rect 428544 339690 428604 340000
rect 430992 339690 431052 340000
rect 428544 339630 428658 339690
rect 418294 337653 418354 339630
rect 415899 337652 415965 337653
rect 415899 337588 415900 337652
rect 415964 337588 415965 337652
rect 415899 337587 415965 337588
rect 418291 337652 418357 337653
rect 418291 337588 418292 337652
rect 418356 337588 418357 337652
rect 418291 337587 418357 337588
rect 414804 308058 414986 308294
rect 415222 308058 415404 308294
rect 414804 272294 415404 308058
rect 414804 272058 414986 272294
rect 415222 272058 415404 272294
rect 414804 236294 415404 272058
rect 414804 236058 414986 236294
rect 415222 236058 415404 236294
rect 414804 200294 415404 236058
rect 414804 200058 414986 200294
rect 415222 200058 415404 200294
rect 414804 164294 415404 200058
rect 414804 164058 414986 164294
rect 415222 164058 415404 164294
rect 414804 128294 415404 164058
rect 414804 128058 414986 128294
rect 415222 128058 415404 128294
rect 414804 92294 415404 128058
rect 414804 92058 414986 92294
rect 415222 92058 415404 92294
rect 414804 56294 415404 92058
rect 414804 56058 414986 56294
rect 415222 56058 415404 56294
rect 414804 20294 415404 56058
rect 414804 20058 414986 20294
rect 415222 20058 415404 20294
rect 414804 -1306 415404 20058
rect 414804 -1542 414986 -1306
rect 415222 -1542 415404 -1306
rect 414804 -1626 415404 -1542
rect 414804 -1862 414986 -1626
rect 415222 -1862 415404 -1626
rect 414804 -1894 415404 -1862
rect 418504 311994 419104 338000
rect 420870 337653 420930 339630
rect 420867 337652 420933 337653
rect 420867 337588 420868 337652
rect 420932 337588 420933 337652
rect 420867 337587 420933 337588
rect 418504 311758 418686 311994
rect 418922 311758 419104 311994
rect 418504 275994 419104 311758
rect 418504 275758 418686 275994
rect 418922 275758 419104 275994
rect 418504 239994 419104 275758
rect 418504 239758 418686 239994
rect 418922 239758 419104 239994
rect 418504 203994 419104 239758
rect 418504 203758 418686 203994
rect 418922 203758 419104 203994
rect 418504 167994 419104 203758
rect 418504 167758 418686 167994
rect 418922 167758 419104 167994
rect 418504 131994 419104 167758
rect 418504 131758 418686 131994
rect 418922 131758 419104 131994
rect 418504 95994 419104 131758
rect 418504 95758 418686 95994
rect 418922 95758 419104 95994
rect 418504 59994 419104 95758
rect 418504 59758 418686 59994
rect 418922 59758 419104 59994
rect 418504 23994 419104 59758
rect 418504 23758 418686 23994
rect 418922 23758 419104 23994
rect 418504 -3226 419104 23758
rect 418504 -3462 418686 -3226
rect 418922 -3462 419104 -3226
rect 418504 -3546 419104 -3462
rect 418504 -3782 418686 -3546
rect 418922 -3782 419104 -3546
rect 418504 -3814 419104 -3782
rect 422204 315694 422804 338000
rect 423446 337381 423506 339630
rect 423443 337380 423509 337381
rect 423443 337316 423444 337380
rect 423508 337316 423509 337380
rect 423443 337315 423509 337316
rect 425654 336973 425714 339630
rect 425651 336972 425717 336973
rect 425651 336908 425652 336972
rect 425716 336908 425717 336972
rect 425651 336907 425717 336908
rect 422204 315458 422386 315694
rect 422622 315458 422804 315694
rect 422204 279694 422804 315458
rect 422204 279458 422386 279694
rect 422622 279458 422804 279694
rect 422204 243694 422804 279458
rect 422204 243458 422386 243694
rect 422622 243458 422804 243694
rect 422204 207694 422804 243458
rect 422204 207458 422386 207694
rect 422622 207458 422804 207694
rect 422204 171694 422804 207458
rect 422204 171458 422386 171694
rect 422622 171458 422804 171694
rect 422204 135694 422804 171458
rect 422204 135458 422386 135694
rect 422622 135458 422804 135694
rect 422204 99694 422804 135458
rect 422204 99458 422386 99694
rect 422622 99458 422804 99694
rect 422204 63694 422804 99458
rect 422204 63458 422386 63694
rect 422622 63458 422804 63694
rect 422204 27694 422804 63458
rect 422204 27458 422386 27694
rect 422622 27458 422804 27694
rect 422204 -5146 422804 27458
rect 422204 -5382 422386 -5146
rect 422622 -5382 422804 -5146
rect 422204 -5466 422804 -5382
rect 422204 -5702 422386 -5466
rect 422622 -5702 422804 -5466
rect 422204 -5734 422804 -5702
rect 425904 319394 426504 338000
rect 428598 337653 428658 339630
rect 430990 339630 431052 339690
rect 433440 339690 433500 340000
rect 435888 339690 435948 340000
rect 438472 339690 438532 340000
rect 433440 339630 433626 339690
rect 430990 337653 431050 339630
rect 428595 337652 428661 337653
rect 428595 337588 428596 337652
rect 428660 337588 428661 337652
rect 428595 337587 428661 337588
rect 430987 337652 431053 337653
rect 430987 337588 430988 337652
rect 431052 337588 431053 337652
rect 430987 337587 431053 337588
rect 425904 319158 426086 319394
rect 426322 319158 426504 319394
rect 425904 283394 426504 319158
rect 425904 283158 426086 283394
rect 426322 283158 426504 283394
rect 425904 247394 426504 283158
rect 425904 247158 426086 247394
rect 426322 247158 426504 247394
rect 425904 211394 426504 247158
rect 425904 211158 426086 211394
rect 426322 211158 426504 211394
rect 425904 175394 426504 211158
rect 425904 175158 426086 175394
rect 426322 175158 426504 175394
rect 425904 139394 426504 175158
rect 425904 139158 426086 139394
rect 426322 139158 426504 139394
rect 425904 103394 426504 139158
rect 425904 103158 426086 103394
rect 426322 103158 426504 103394
rect 425904 67394 426504 103158
rect 425904 67158 426086 67394
rect 426322 67158 426504 67394
rect 425904 31394 426504 67158
rect 425904 31158 426086 31394
rect 426322 31158 426504 31394
rect 407904 -6342 408086 -6106
rect 408322 -6342 408504 -6106
rect 407904 -6426 408504 -6342
rect 407904 -6662 408086 -6426
rect 408322 -6662 408504 -6426
rect 407904 -7654 408504 -6662
rect 425904 -7066 426504 31158
rect 432804 326294 433404 338000
rect 433566 337109 433626 339630
rect 435774 339630 435948 339690
rect 438350 339630 438532 339690
rect 440920 339690 440980 340000
rect 443368 339690 443428 340000
rect 445952 339690 446012 340000
rect 440920 339630 440986 339690
rect 435774 337653 435834 339630
rect 435771 337652 435837 337653
rect 435771 337588 435772 337652
rect 435836 337588 435837 337652
rect 435771 337587 435837 337588
rect 433563 337108 433629 337109
rect 433563 337044 433564 337108
rect 433628 337044 433629 337108
rect 433563 337043 433629 337044
rect 432804 326058 432986 326294
rect 433222 326058 433404 326294
rect 432804 290294 433404 326058
rect 432804 290058 432986 290294
rect 433222 290058 433404 290294
rect 432804 254294 433404 290058
rect 432804 254058 432986 254294
rect 433222 254058 433404 254294
rect 432804 218294 433404 254058
rect 432804 218058 432986 218294
rect 433222 218058 433404 218294
rect 432804 182294 433404 218058
rect 432804 182058 432986 182294
rect 433222 182058 433404 182294
rect 432804 146294 433404 182058
rect 432804 146058 432986 146294
rect 433222 146058 433404 146294
rect 432804 110294 433404 146058
rect 432804 110058 432986 110294
rect 433222 110058 433404 110294
rect 432804 74294 433404 110058
rect 432804 74058 432986 74294
rect 433222 74058 433404 74294
rect 432804 38294 433404 74058
rect 432804 38058 432986 38294
rect 433222 38058 433404 38294
rect 432804 2294 433404 38058
rect 432804 2058 432986 2294
rect 433222 2058 433404 2294
rect 432804 -346 433404 2058
rect 432804 -582 432986 -346
rect 433222 -582 433404 -346
rect 432804 -666 433404 -582
rect 432804 -902 432986 -666
rect 433222 -902 433404 -666
rect 432804 -1894 433404 -902
rect 436504 329994 437104 338000
rect 438350 337653 438410 339630
rect 438347 337652 438413 337653
rect 438347 337588 438348 337652
rect 438412 337588 438413 337652
rect 438347 337587 438413 337588
rect 436504 329758 436686 329994
rect 436922 329758 437104 329994
rect 436504 293994 437104 329758
rect 436504 293758 436686 293994
rect 436922 293758 437104 293994
rect 436504 257994 437104 293758
rect 436504 257758 436686 257994
rect 436922 257758 437104 257994
rect 436504 221994 437104 257758
rect 436504 221758 436686 221994
rect 436922 221758 437104 221994
rect 436504 185994 437104 221758
rect 436504 185758 436686 185994
rect 436922 185758 437104 185994
rect 436504 149994 437104 185758
rect 436504 149758 436686 149994
rect 436922 149758 437104 149994
rect 436504 113994 437104 149758
rect 436504 113758 436686 113994
rect 436922 113758 437104 113994
rect 436504 77994 437104 113758
rect 436504 77758 436686 77994
rect 436922 77758 437104 77994
rect 436504 41994 437104 77758
rect 436504 41758 436686 41994
rect 436922 41758 437104 41994
rect 436504 5994 437104 41758
rect 436504 5758 436686 5994
rect 436922 5758 437104 5994
rect 436504 -2266 437104 5758
rect 436504 -2502 436686 -2266
rect 436922 -2502 437104 -2266
rect 436504 -2586 437104 -2502
rect 436504 -2822 436686 -2586
rect 436922 -2822 437104 -2586
rect 436504 -3814 437104 -2822
rect 440204 333694 440804 338000
rect 440926 337109 440986 339630
rect 443318 339630 443428 339690
rect 445894 339630 446012 339690
rect 443318 337245 443378 339630
rect 443904 337394 444504 338000
rect 445894 337653 445954 339630
rect 445891 337652 445957 337653
rect 445891 337588 445892 337652
rect 445956 337588 445957 337652
rect 445891 337587 445957 337588
rect 443315 337244 443381 337245
rect 443315 337180 443316 337244
rect 443380 337180 443381 337244
rect 443315 337179 443381 337180
rect 443904 337158 444086 337394
rect 444322 337158 444504 337394
rect 440923 337108 440989 337109
rect 440923 337044 440924 337108
rect 440988 337044 440989 337108
rect 440923 337043 440989 337044
rect 440204 333458 440386 333694
rect 440622 333458 440804 333694
rect 440204 297694 440804 333458
rect 440204 297458 440386 297694
rect 440622 297458 440804 297694
rect 440204 261694 440804 297458
rect 440204 261458 440386 261694
rect 440622 261458 440804 261694
rect 440204 225694 440804 261458
rect 440204 225458 440386 225694
rect 440622 225458 440804 225694
rect 440204 189694 440804 225458
rect 440204 189458 440386 189694
rect 440622 189458 440804 189694
rect 440204 153694 440804 189458
rect 440204 153458 440386 153694
rect 440622 153458 440804 153694
rect 440204 117694 440804 153458
rect 440204 117458 440386 117694
rect 440622 117458 440804 117694
rect 440204 81694 440804 117458
rect 440204 81458 440386 81694
rect 440622 81458 440804 81694
rect 440204 45694 440804 81458
rect 440204 45458 440386 45694
rect 440622 45458 440804 45694
rect 440204 9694 440804 45458
rect 440204 9458 440386 9694
rect 440622 9458 440804 9694
rect 440204 -4186 440804 9458
rect 440204 -4422 440386 -4186
rect 440622 -4422 440804 -4186
rect 440204 -4506 440804 -4422
rect 440204 -4742 440386 -4506
rect 440622 -4742 440804 -4506
rect 440204 -5734 440804 -4742
rect 443904 301394 444504 337158
rect 443904 301158 444086 301394
rect 444322 301158 444504 301394
rect 443904 265394 444504 301158
rect 443904 265158 444086 265394
rect 444322 265158 444504 265394
rect 443904 229394 444504 265158
rect 443904 229158 444086 229394
rect 444322 229158 444504 229394
rect 443904 193394 444504 229158
rect 443904 193158 444086 193394
rect 444322 193158 444504 193394
rect 443904 157394 444504 193158
rect 443904 157158 444086 157394
rect 444322 157158 444504 157394
rect 443904 121394 444504 157158
rect 443904 121158 444086 121394
rect 444322 121158 444504 121394
rect 443904 85394 444504 121158
rect 443904 85158 444086 85394
rect 444322 85158 444504 85394
rect 443904 49394 444504 85158
rect 443904 49158 444086 49394
rect 444322 49158 444504 49394
rect 443904 13394 444504 49158
rect 443904 13158 444086 13394
rect 444322 13158 444504 13394
rect 425904 -7302 426086 -7066
rect 426322 -7302 426504 -7066
rect 425904 -7386 426504 -7302
rect 425904 -7622 426086 -7386
rect 426322 -7622 426504 -7386
rect 425904 -7654 426504 -7622
rect 443904 -6106 444504 13158
rect 450804 308294 451404 338000
rect 450804 308058 450986 308294
rect 451222 308058 451404 308294
rect 450804 272294 451404 308058
rect 450804 272058 450986 272294
rect 451222 272058 451404 272294
rect 450804 236294 451404 272058
rect 450804 236058 450986 236294
rect 451222 236058 451404 236294
rect 450804 200294 451404 236058
rect 450804 200058 450986 200294
rect 451222 200058 451404 200294
rect 450804 164294 451404 200058
rect 450804 164058 450986 164294
rect 451222 164058 451404 164294
rect 450804 128294 451404 164058
rect 450804 128058 450986 128294
rect 451222 128058 451404 128294
rect 450804 92294 451404 128058
rect 450804 92058 450986 92294
rect 451222 92058 451404 92294
rect 450804 56294 451404 92058
rect 450804 56058 450986 56294
rect 451222 56058 451404 56294
rect 450804 20294 451404 56058
rect 450804 20058 450986 20294
rect 451222 20058 451404 20294
rect 450804 -1306 451404 20058
rect 450804 -1542 450986 -1306
rect 451222 -1542 451404 -1306
rect 450804 -1626 451404 -1542
rect 450804 -1862 450986 -1626
rect 451222 -1862 451404 -1626
rect 450804 -1894 451404 -1862
rect 454504 311994 455104 338000
rect 454504 311758 454686 311994
rect 454922 311758 455104 311994
rect 454504 275994 455104 311758
rect 454504 275758 454686 275994
rect 454922 275758 455104 275994
rect 454504 239994 455104 275758
rect 454504 239758 454686 239994
rect 454922 239758 455104 239994
rect 454504 203994 455104 239758
rect 454504 203758 454686 203994
rect 454922 203758 455104 203994
rect 454504 167994 455104 203758
rect 454504 167758 454686 167994
rect 454922 167758 455104 167994
rect 454504 131994 455104 167758
rect 454504 131758 454686 131994
rect 454922 131758 455104 131994
rect 454504 95994 455104 131758
rect 454504 95758 454686 95994
rect 454922 95758 455104 95994
rect 454504 59994 455104 95758
rect 454504 59758 454686 59994
rect 454922 59758 455104 59994
rect 454504 23994 455104 59758
rect 454504 23758 454686 23994
rect 454922 23758 455104 23994
rect 454504 -3226 455104 23758
rect 454504 -3462 454686 -3226
rect 454922 -3462 455104 -3226
rect 454504 -3546 455104 -3462
rect 454504 -3782 454686 -3546
rect 454922 -3782 455104 -3546
rect 454504 -3814 455104 -3782
rect 458204 315694 458804 338000
rect 458204 315458 458386 315694
rect 458622 315458 458804 315694
rect 458204 279694 458804 315458
rect 458204 279458 458386 279694
rect 458622 279458 458804 279694
rect 458204 243694 458804 279458
rect 458204 243458 458386 243694
rect 458622 243458 458804 243694
rect 458204 207694 458804 243458
rect 458204 207458 458386 207694
rect 458622 207458 458804 207694
rect 458204 171694 458804 207458
rect 458204 171458 458386 171694
rect 458622 171458 458804 171694
rect 458204 135694 458804 171458
rect 458204 135458 458386 135694
rect 458622 135458 458804 135694
rect 458204 99694 458804 135458
rect 458204 99458 458386 99694
rect 458622 99458 458804 99694
rect 458204 63694 458804 99458
rect 458204 63458 458386 63694
rect 458622 63458 458804 63694
rect 458204 27694 458804 63458
rect 458204 27458 458386 27694
rect 458622 27458 458804 27694
rect 458204 -5146 458804 27458
rect 458204 -5382 458386 -5146
rect 458622 -5382 458804 -5146
rect 458204 -5466 458804 -5382
rect 458204 -5702 458386 -5466
rect 458622 -5702 458804 -5466
rect 458204 -5734 458804 -5702
rect 461904 319394 462504 338000
rect 461904 319158 462086 319394
rect 462322 319158 462504 319394
rect 461904 283394 462504 319158
rect 461904 283158 462086 283394
rect 462322 283158 462504 283394
rect 461904 247394 462504 283158
rect 461904 247158 462086 247394
rect 462322 247158 462504 247394
rect 461904 211394 462504 247158
rect 461904 211158 462086 211394
rect 462322 211158 462504 211394
rect 461904 175394 462504 211158
rect 461904 175158 462086 175394
rect 462322 175158 462504 175394
rect 461904 139394 462504 175158
rect 461904 139158 462086 139394
rect 462322 139158 462504 139394
rect 461904 103394 462504 139158
rect 461904 103158 462086 103394
rect 462322 103158 462504 103394
rect 461904 67394 462504 103158
rect 461904 67158 462086 67394
rect 462322 67158 462504 67394
rect 461904 31394 462504 67158
rect 461904 31158 462086 31394
rect 462322 31158 462504 31394
rect 443904 -6342 444086 -6106
rect 444322 -6342 444504 -6106
rect 443904 -6426 444504 -6342
rect 443904 -6662 444086 -6426
rect 444322 -6662 444504 -6426
rect 443904 -7654 444504 -6662
rect 461904 -7066 462504 31158
rect 468804 326294 469404 338000
rect 468804 326058 468986 326294
rect 469222 326058 469404 326294
rect 468804 290294 469404 326058
rect 468804 290058 468986 290294
rect 469222 290058 469404 290294
rect 468804 254294 469404 290058
rect 468804 254058 468986 254294
rect 469222 254058 469404 254294
rect 468804 218294 469404 254058
rect 468804 218058 468986 218294
rect 469222 218058 469404 218294
rect 468804 182294 469404 218058
rect 468804 182058 468986 182294
rect 469222 182058 469404 182294
rect 468804 146294 469404 182058
rect 468804 146058 468986 146294
rect 469222 146058 469404 146294
rect 468804 110294 469404 146058
rect 468804 110058 468986 110294
rect 469222 110058 469404 110294
rect 468804 74294 469404 110058
rect 468804 74058 468986 74294
rect 469222 74058 469404 74294
rect 468804 38294 469404 74058
rect 468804 38058 468986 38294
rect 469222 38058 469404 38294
rect 468804 2294 469404 38058
rect 468804 2058 468986 2294
rect 469222 2058 469404 2294
rect 468804 -346 469404 2058
rect 468804 -582 468986 -346
rect 469222 -582 469404 -346
rect 468804 -666 469404 -582
rect 468804 -902 468986 -666
rect 469222 -902 469404 -666
rect 468804 -1894 469404 -902
rect 472504 329994 473104 338000
rect 472504 329758 472686 329994
rect 472922 329758 473104 329994
rect 472504 293994 473104 329758
rect 472504 293758 472686 293994
rect 472922 293758 473104 293994
rect 472504 257994 473104 293758
rect 472504 257758 472686 257994
rect 472922 257758 473104 257994
rect 472504 221994 473104 257758
rect 472504 221758 472686 221994
rect 472922 221758 473104 221994
rect 472504 185994 473104 221758
rect 472504 185758 472686 185994
rect 472922 185758 473104 185994
rect 472504 149994 473104 185758
rect 472504 149758 472686 149994
rect 472922 149758 473104 149994
rect 472504 113994 473104 149758
rect 472504 113758 472686 113994
rect 472922 113758 473104 113994
rect 472504 77994 473104 113758
rect 472504 77758 472686 77994
rect 472922 77758 473104 77994
rect 472504 41994 473104 77758
rect 472504 41758 472686 41994
rect 472922 41758 473104 41994
rect 472504 5994 473104 41758
rect 472504 5758 472686 5994
rect 472922 5758 473104 5994
rect 472504 -2266 473104 5758
rect 472504 -2502 472686 -2266
rect 472922 -2502 473104 -2266
rect 472504 -2586 473104 -2502
rect 472504 -2822 472686 -2586
rect 472922 -2822 473104 -2586
rect 472504 -3814 473104 -2822
rect 476204 333694 476804 338000
rect 476204 333458 476386 333694
rect 476622 333458 476804 333694
rect 476204 297694 476804 333458
rect 476204 297458 476386 297694
rect 476622 297458 476804 297694
rect 476204 261694 476804 297458
rect 476204 261458 476386 261694
rect 476622 261458 476804 261694
rect 476204 225694 476804 261458
rect 476204 225458 476386 225694
rect 476622 225458 476804 225694
rect 476204 189694 476804 225458
rect 476204 189458 476386 189694
rect 476622 189458 476804 189694
rect 476204 153694 476804 189458
rect 476204 153458 476386 153694
rect 476622 153458 476804 153694
rect 476204 117694 476804 153458
rect 476204 117458 476386 117694
rect 476622 117458 476804 117694
rect 476204 81694 476804 117458
rect 476204 81458 476386 81694
rect 476622 81458 476804 81694
rect 476204 45694 476804 81458
rect 476204 45458 476386 45694
rect 476622 45458 476804 45694
rect 476204 9694 476804 45458
rect 476204 9458 476386 9694
rect 476622 9458 476804 9694
rect 476204 -4186 476804 9458
rect 476204 -4422 476386 -4186
rect 476622 -4422 476804 -4186
rect 476204 -4506 476804 -4422
rect 476204 -4742 476386 -4506
rect 476622 -4742 476804 -4506
rect 476204 -5734 476804 -4742
rect 479904 337394 480504 373158
rect 479904 337158 480086 337394
rect 480322 337158 480504 337394
rect 479904 301394 480504 337158
rect 479904 301158 480086 301394
rect 480322 301158 480504 301394
rect 479904 265394 480504 301158
rect 479904 265158 480086 265394
rect 480322 265158 480504 265394
rect 479904 229394 480504 265158
rect 479904 229158 480086 229394
rect 480322 229158 480504 229394
rect 479904 193394 480504 229158
rect 479904 193158 480086 193394
rect 480322 193158 480504 193394
rect 479904 157394 480504 193158
rect 479904 157158 480086 157394
rect 480322 157158 480504 157394
rect 479904 121394 480504 157158
rect 479904 121158 480086 121394
rect 480322 121158 480504 121394
rect 479904 85394 480504 121158
rect 479904 85158 480086 85394
rect 480322 85158 480504 85394
rect 479904 49394 480504 85158
rect 479904 49158 480086 49394
rect 480322 49158 480504 49394
rect 479904 13394 480504 49158
rect 479904 13158 480086 13394
rect 480322 13158 480504 13394
rect 461904 -7302 462086 -7066
rect 462322 -7302 462504 -7066
rect 461904 -7386 462504 -7302
rect 461904 -7622 462086 -7386
rect 462322 -7622 462504 -7386
rect 461904 -7654 462504 -7622
rect 479904 -6106 480504 13158
rect 486804 705798 487404 705830
rect 486804 705562 486986 705798
rect 487222 705562 487404 705798
rect 486804 705478 487404 705562
rect 486804 705242 486986 705478
rect 487222 705242 487404 705478
rect 486804 668294 487404 705242
rect 486804 668058 486986 668294
rect 487222 668058 487404 668294
rect 486804 632294 487404 668058
rect 486804 632058 486986 632294
rect 487222 632058 487404 632294
rect 486804 596294 487404 632058
rect 486804 596058 486986 596294
rect 487222 596058 487404 596294
rect 486804 560294 487404 596058
rect 486804 560058 486986 560294
rect 487222 560058 487404 560294
rect 486804 524294 487404 560058
rect 486804 524058 486986 524294
rect 487222 524058 487404 524294
rect 486804 488294 487404 524058
rect 486804 488058 486986 488294
rect 487222 488058 487404 488294
rect 486804 452294 487404 488058
rect 486804 452058 486986 452294
rect 487222 452058 487404 452294
rect 486804 416294 487404 452058
rect 486804 416058 486986 416294
rect 487222 416058 487404 416294
rect 486804 380294 487404 416058
rect 486804 380058 486986 380294
rect 487222 380058 487404 380294
rect 486804 344294 487404 380058
rect 486804 344058 486986 344294
rect 487222 344058 487404 344294
rect 486804 308294 487404 344058
rect 486804 308058 486986 308294
rect 487222 308058 487404 308294
rect 486804 272294 487404 308058
rect 486804 272058 486986 272294
rect 487222 272058 487404 272294
rect 486804 236294 487404 272058
rect 486804 236058 486986 236294
rect 487222 236058 487404 236294
rect 486804 200294 487404 236058
rect 486804 200058 486986 200294
rect 487222 200058 487404 200294
rect 486804 164294 487404 200058
rect 486804 164058 486986 164294
rect 487222 164058 487404 164294
rect 486804 128294 487404 164058
rect 486804 128058 486986 128294
rect 487222 128058 487404 128294
rect 486804 92294 487404 128058
rect 486804 92058 486986 92294
rect 487222 92058 487404 92294
rect 486804 56294 487404 92058
rect 486804 56058 486986 56294
rect 487222 56058 487404 56294
rect 486804 20294 487404 56058
rect 486804 20058 486986 20294
rect 487222 20058 487404 20294
rect 486804 -1306 487404 20058
rect 486804 -1542 486986 -1306
rect 487222 -1542 487404 -1306
rect 486804 -1626 487404 -1542
rect 486804 -1862 486986 -1626
rect 487222 -1862 487404 -1626
rect 486804 -1894 487404 -1862
rect 490504 671994 491104 707162
rect 490504 671758 490686 671994
rect 490922 671758 491104 671994
rect 490504 635994 491104 671758
rect 490504 635758 490686 635994
rect 490922 635758 491104 635994
rect 490504 599994 491104 635758
rect 490504 599758 490686 599994
rect 490922 599758 491104 599994
rect 490504 563994 491104 599758
rect 490504 563758 490686 563994
rect 490922 563758 491104 563994
rect 490504 527994 491104 563758
rect 490504 527758 490686 527994
rect 490922 527758 491104 527994
rect 490504 491994 491104 527758
rect 490504 491758 490686 491994
rect 490922 491758 491104 491994
rect 490504 455994 491104 491758
rect 490504 455758 490686 455994
rect 490922 455758 491104 455994
rect 490504 419994 491104 455758
rect 490504 419758 490686 419994
rect 490922 419758 491104 419994
rect 490504 383994 491104 419758
rect 490504 383758 490686 383994
rect 490922 383758 491104 383994
rect 490504 347994 491104 383758
rect 490504 347758 490686 347994
rect 490922 347758 491104 347994
rect 490504 311994 491104 347758
rect 490504 311758 490686 311994
rect 490922 311758 491104 311994
rect 490504 275994 491104 311758
rect 490504 275758 490686 275994
rect 490922 275758 491104 275994
rect 490504 239994 491104 275758
rect 490504 239758 490686 239994
rect 490922 239758 491104 239994
rect 490504 203994 491104 239758
rect 490504 203758 490686 203994
rect 490922 203758 491104 203994
rect 490504 167994 491104 203758
rect 490504 167758 490686 167994
rect 490922 167758 491104 167994
rect 490504 131994 491104 167758
rect 490504 131758 490686 131994
rect 490922 131758 491104 131994
rect 490504 95994 491104 131758
rect 490504 95758 490686 95994
rect 490922 95758 491104 95994
rect 490504 59994 491104 95758
rect 490504 59758 490686 59994
rect 490922 59758 491104 59994
rect 490504 23994 491104 59758
rect 490504 23758 490686 23994
rect 490922 23758 491104 23994
rect 490504 -3226 491104 23758
rect 490504 -3462 490686 -3226
rect 490922 -3462 491104 -3226
rect 490504 -3546 491104 -3462
rect 490504 -3782 490686 -3546
rect 490922 -3782 491104 -3546
rect 490504 -3814 491104 -3782
rect 494204 675694 494804 709082
rect 494204 675458 494386 675694
rect 494622 675458 494804 675694
rect 494204 639694 494804 675458
rect 494204 639458 494386 639694
rect 494622 639458 494804 639694
rect 494204 603694 494804 639458
rect 494204 603458 494386 603694
rect 494622 603458 494804 603694
rect 494204 567694 494804 603458
rect 494204 567458 494386 567694
rect 494622 567458 494804 567694
rect 494204 531694 494804 567458
rect 494204 531458 494386 531694
rect 494622 531458 494804 531694
rect 494204 495694 494804 531458
rect 494204 495458 494386 495694
rect 494622 495458 494804 495694
rect 494204 459694 494804 495458
rect 494204 459458 494386 459694
rect 494622 459458 494804 459694
rect 494204 423694 494804 459458
rect 494204 423458 494386 423694
rect 494622 423458 494804 423694
rect 494204 387694 494804 423458
rect 494204 387458 494386 387694
rect 494622 387458 494804 387694
rect 494204 351694 494804 387458
rect 494204 351458 494386 351694
rect 494622 351458 494804 351694
rect 494204 315694 494804 351458
rect 494204 315458 494386 315694
rect 494622 315458 494804 315694
rect 494204 279694 494804 315458
rect 494204 279458 494386 279694
rect 494622 279458 494804 279694
rect 494204 243694 494804 279458
rect 494204 243458 494386 243694
rect 494622 243458 494804 243694
rect 494204 207694 494804 243458
rect 494204 207458 494386 207694
rect 494622 207458 494804 207694
rect 494204 171694 494804 207458
rect 494204 171458 494386 171694
rect 494622 171458 494804 171694
rect 494204 135694 494804 171458
rect 494204 135458 494386 135694
rect 494622 135458 494804 135694
rect 494204 99694 494804 135458
rect 494204 99458 494386 99694
rect 494622 99458 494804 99694
rect 494204 63694 494804 99458
rect 494204 63458 494386 63694
rect 494622 63458 494804 63694
rect 494204 27694 494804 63458
rect 494204 27458 494386 27694
rect 494622 27458 494804 27694
rect 494204 -5146 494804 27458
rect 494204 -5382 494386 -5146
rect 494622 -5382 494804 -5146
rect 494204 -5466 494804 -5382
rect 494204 -5702 494386 -5466
rect 494622 -5702 494804 -5466
rect 494204 -5734 494804 -5702
rect 497904 679394 498504 711002
rect 515904 710598 516504 711590
rect 515904 710362 516086 710598
rect 516322 710362 516504 710598
rect 515904 710278 516504 710362
rect 515904 710042 516086 710278
rect 516322 710042 516504 710278
rect 512204 708678 512804 709670
rect 512204 708442 512386 708678
rect 512622 708442 512804 708678
rect 512204 708358 512804 708442
rect 512204 708122 512386 708358
rect 512622 708122 512804 708358
rect 508504 706758 509104 707750
rect 508504 706522 508686 706758
rect 508922 706522 509104 706758
rect 508504 706438 509104 706522
rect 508504 706202 508686 706438
rect 508922 706202 509104 706438
rect 497904 679158 498086 679394
rect 498322 679158 498504 679394
rect 497904 643394 498504 679158
rect 497904 643158 498086 643394
rect 498322 643158 498504 643394
rect 497904 607394 498504 643158
rect 497904 607158 498086 607394
rect 498322 607158 498504 607394
rect 497904 571394 498504 607158
rect 497904 571158 498086 571394
rect 498322 571158 498504 571394
rect 497904 535394 498504 571158
rect 497904 535158 498086 535394
rect 498322 535158 498504 535394
rect 497904 499394 498504 535158
rect 497904 499158 498086 499394
rect 498322 499158 498504 499394
rect 497904 463394 498504 499158
rect 497904 463158 498086 463394
rect 498322 463158 498504 463394
rect 497904 427394 498504 463158
rect 497904 427158 498086 427394
rect 498322 427158 498504 427394
rect 497904 391394 498504 427158
rect 497904 391158 498086 391394
rect 498322 391158 498504 391394
rect 497904 355394 498504 391158
rect 497904 355158 498086 355394
rect 498322 355158 498504 355394
rect 497904 319394 498504 355158
rect 497904 319158 498086 319394
rect 498322 319158 498504 319394
rect 497904 283394 498504 319158
rect 497904 283158 498086 283394
rect 498322 283158 498504 283394
rect 497904 247394 498504 283158
rect 497904 247158 498086 247394
rect 498322 247158 498504 247394
rect 497904 211394 498504 247158
rect 497904 211158 498086 211394
rect 498322 211158 498504 211394
rect 497904 175394 498504 211158
rect 497904 175158 498086 175394
rect 498322 175158 498504 175394
rect 497904 139394 498504 175158
rect 497904 139158 498086 139394
rect 498322 139158 498504 139394
rect 497904 103394 498504 139158
rect 497904 103158 498086 103394
rect 498322 103158 498504 103394
rect 497904 67394 498504 103158
rect 497904 67158 498086 67394
rect 498322 67158 498504 67394
rect 497904 31394 498504 67158
rect 497904 31158 498086 31394
rect 498322 31158 498504 31394
rect 479904 -6342 480086 -6106
rect 480322 -6342 480504 -6106
rect 479904 -6426 480504 -6342
rect 479904 -6662 480086 -6426
rect 480322 -6662 480504 -6426
rect 479904 -7654 480504 -6662
rect 497904 -7066 498504 31158
rect 504804 704838 505404 705830
rect 504804 704602 504986 704838
rect 505222 704602 505404 704838
rect 504804 704518 505404 704602
rect 504804 704282 504986 704518
rect 505222 704282 505404 704518
rect 504804 686294 505404 704282
rect 504804 686058 504986 686294
rect 505222 686058 505404 686294
rect 504804 650294 505404 686058
rect 504804 650058 504986 650294
rect 505222 650058 505404 650294
rect 504804 614294 505404 650058
rect 504804 614058 504986 614294
rect 505222 614058 505404 614294
rect 504804 578294 505404 614058
rect 504804 578058 504986 578294
rect 505222 578058 505404 578294
rect 504804 542294 505404 578058
rect 504804 542058 504986 542294
rect 505222 542058 505404 542294
rect 504804 506294 505404 542058
rect 504804 506058 504986 506294
rect 505222 506058 505404 506294
rect 504804 470294 505404 506058
rect 504804 470058 504986 470294
rect 505222 470058 505404 470294
rect 504804 434294 505404 470058
rect 504804 434058 504986 434294
rect 505222 434058 505404 434294
rect 504804 398294 505404 434058
rect 504804 398058 504986 398294
rect 505222 398058 505404 398294
rect 504804 362294 505404 398058
rect 504804 362058 504986 362294
rect 505222 362058 505404 362294
rect 504804 326294 505404 362058
rect 504804 326058 504986 326294
rect 505222 326058 505404 326294
rect 504804 290294 505404 326058
rect 504804 290058 504986 290294
rect 505222 290058 505404 290294
rect 504804 254294 505404 290058
rect 504804 254058 504986 254294
rect 505222 254058 505404 254294
rect 504804 218294 505404 254058
rect 504804 218058 504986 218294
rect 505222 218058 505404 218294
rect 504804 182294 505404 218058
rect 504804 182058 504986 182294
rect 505222 182058 505404 182294
rect 504804 146294 505404 182058
rect 504804 146058 504986 146294
rect 505222 146058 505404 146294
rect 504804 110294 505404 146058
rect 504804 110058 504986 110294
rect 505222 110058 505404 110294
rect 504804 74294 505404 110058
rect 504804 74058 504986 74294
rect 505222 74058 505404 74294
rect 504804 38294 505404 74058
rect 504804 38058 504986 38294
rect 505222 38058 505404 38294
rect 504804 2294 505404 38058
rect 504804 2058 504986 2294
rect 505222 2058 505404 2294
rect 504804 -346 505404 2058
rect 504804 -582 504986 -346
rect 505222 -582 505404 -346
rect 504804 -666 505404 -582
rect 504804 -902 504986 -666
rect 505222 -902 505404 -666
rect 504804 -1894 505404 -902
rect 508504 689994 509104 706202
rect 508504 689758 508686 689994
rect 508922 689758 509104 689994
rect 508504 653994 509104 689758
rect 508504 653758 508686 653994
rect 508922 653758 509104 653994
rect 508504 617994 509104 653758
rect 508504 617758 508686 617994
rect 508922 617758 509104 617994
rect 508504 581994 509104 617758
rect 508504 581758 508686 581994
rect 508922 581758 509104 581994
rect 508504 545994 509104 581758
rect 508504 545758 508686 545994
rect 508922 545758 509104 545994
rect 508504 509994 509104 545758
rect 508504 509758 508686 509994
rect 508922 509758 509104 509994
rect 508504 473994 509104 509758
rect 508504 473758 508686 473994
rect 508922 473758 509104 473994
rect 508504 437994 509104 473758
rect 508504 437758 508686 437994
rect 508922 437758 509104 437994
rect 508504 401994 509104 437758
rect 508504 401758 508686 401994
rect 508922 401758 509104 401994
rect 508504 365994 509104 401758
rect 508504 365758 508686 365994
rect 508922 365758 509104 365994
rect 508504 329994 509104 365758
rect 508504 329758 508686 329994
rect 508922 329758 509104 329994
rect 508504 293994 509104 329758
rect 508504 293758 508686 293994
rect 508922 293758 509104 293994
rect 508504 257994 509104 293758
rect 508504 257758 508686 257994
rect 508922 257758 509104 257994
rect 508504 221994 509104 257758
rect 508504 221758 508686 221994
rect 508922 221758 509104 221994
rect 508504 185994 509104 221758
rect 508504 185758 508686 185994
rect 508922 185758 509104 185994
rect 508504 149994 509104 185758
rect 508504 149758 508686 149994
rect 508922 149758 509104 149994
rect 508504 113994 509104 149758
rect 508504 113758 508686 113994
rect 508922 113758 509104 113994
rect 508504 77994 509104 113758
rect 508504 77758 508686 77994
rect 508922 77758 509104 77994
rect 508504 41994 509104 77758
rect 508504 41758 508686 41994
rect 508922 41758 509104 41994
rect 508504 5994 509104 41758
rect 508504 5758 508686 5994
rect 508922 5758 509104 5994
rect 508504 -2266 509104 5758
rect 508504 -2502 508686 -2266
rect 508922 -2502 509104 -2266
rect 508504 -2586 509104 -2502
rect 508504 -2822 508686 -2586
rect 508922 -2822 509104 -2586
rect 508504 -3814 509104 -2822
rect 512204 693694 512804 708122
rect 512204 693458 512386 693694
rect 512622 693458 512804 693694
rect 512204 657694 512804 693458
rect 512204 657458 512386 657694
rect 512622 657458 512804 657694
rect 512204 621694 512804 657458
rect 512204 621458 512386 621694
rect 512622 621458 512804 621694
rect 512204 585694 512804 621458
rect 512204 585458 512386 585694
rect 512622 585458 512804 585694
rect 512204 549694 512804 585458
rect 512204 549458 512386 549694
rect 512622 549458 512804 549694
rect 512204 513694 512804 549458
rect 512204 513458 512386 513694
rect 512622 513458 512804 513694
rect 512204 477694 512804 513458
rect 512204 477458 512386 477694
rect 512622 477458 512804 477694
rect 512204 441694 512804 477458
rect 512204 441458 512386 441694
rect 512622 441458 512804 441694
rect 512204 405694 512804 441458
rect 512204 405458 512386 405694
rect 512622 405458 512804 405694
rect 512204 369694 512804 405458
rect 512204 369458 512386 369694
rect 512622 369458 512804 369694
rect 512204 333694 512804 369458
rect 512204 333458 512386 333694
rect 512622 333458 512804 333694
rect 512204 297694 512804 333458
rect 512204 297458 512386 297694
rect 512622 297458 512804 297694
rect 512204 261694 512804 297458
rect 512204 261458 512386 261694
rect 512622 261458 512804 261694
rect 512204 225694 512804 261458
rect 512204 225458 512386 225694
rect 512622 225458 512804 225694
rect 512204 189694 512804 225458
rect 512204 189458 512386 189694
rect 512622 189458 512804 189694
rect 512204 153694 512804 189458
rect 512204 153458 512386 153694
rect 512622 153458 512804 153694
rect 512204 117694 512804 153458
rect 512204 117458 512386 117694
rect 512622 117458 512804 117694
rect 512204 81694 512804 117458
rect 512204 81458 512386 81694
rect 512622 81458 512804 81694
rect 512204 45694 512804 81458
rect 512204 45458 512386 45694
rect 512622 45458 512804 45694
rect 512204 9694 512804 45458
rect 512204 9458 512386 9694
rect 512622 9458 512804 9694
rect 512204 -4186 512804 9458
rect 512204 -4422 512386 -4186
rect 512622 -4422 512804 -4186
rect 512204 -4506 512804 -4422
rect 512204 -4742 512386 -4506
rect 512622 -4742 512804 -4506
rect 512204 -5734 512804 -4742
rect 515904 697394 516504 710042
rect 533904 711558 534504 711590
rect 533904 711322 534086 711558
rect 534322 711322 534504 711558
rect 533904 711238 534504 711322
rect 533904 711002 534086 711238
rect 534322 711002 534504 711238
rect 530204 709638 530804 709670
rect 530204 709402 530386 709638
rect 530622 709402 530804 709638
rect 530204 709318 530804 709402
rect 530204 709082 530386 709318
rect 530622 709082 530804 709318
rect 526504 707718 527104 707750
rect 526504 707482 526686 707718
rect 526922 707482 527104 707718
rect 526504 707398 527104 707482
rect 526504 707162 526686 707398
rect 526922 707162 527104 707398
rect 515904 697158 516086 697394
rect 516322 697158 516504 697394
rect 515904 661394 516504 697158
rect 515904 661158 516086 661394
rect 516322 661158 516504 661394
rect 515904 625394 516504 661158
rect 515904 625158 516086 625394
rect 516322 625158 516504 625394
rect 515904 589394 516504 625158
rect 515904 589158 516086 589394
rect 516322 589158 516504 589394
rect 515904 553394 516504 589158
rect 515904 553158 516086 553394
rect 516322 553158 516504 553394
rect 515904 517394 516504 553158
rect 515904 517158 516086 517394
rect 516322 517158 516504 517394
rect 515904 481394 516504 517158
rect 515904 481158 516086 481394
rect 516322 481158 516504 481394
rect 515904 445394 516504 481158
rect 515904 445158 516086 445394
rect 516322 445158 516504 445394
rect 515904 409394 516504 445158
rect 515904 409158 516086 409394
rect 516322 409158 516504 409394
rect 515904 373394 516504 409158
rect 515904 373158 516086 373394
rect 516322 373158 516504 373394
rect 515904 337394 516504 373158
rect 515904 337158 516086 337394
rect 516322 337158 516504 337394
rect 515904 301394 516504 337158
rect 515904 301158 516086 301394
rect 516322 301158 516504 301394
rect 515904 265394 516504 301158
rect 515904 265158 516086 265394
rect 516322 265158 516504 265394
rect 515904 229394 516504 265158
rect 515904 229158 516086 229394
rect 516322 229158 516504 229394
rect 515904 193394 516504 229158
rect 515904 193158 516086 193394
rect 516322 193158 516504 193394
rect 515904 157394 516504 193158
rect 515904 157158 516086 157394
rect 516322 157158 516504 157394
rect 515904 121394 516504 157158
rect 515904 121158 516086 121394
rect 516322 121158 516504 121394
rect 515904 85394 516504 121158
rect 515904 85158 516086 85394
rect 516322 85158 516504 85394
rect 515904 49394 516504 85158
rect 515904 49158 516086 49394
rect 516322 49158 516504 49394
rect 515904 13394 516504 49158
rect 515904 13158 516086 13394
rect 516322 13158 516504 13394
rect 497904 -7302 498086 -7066
rect 498322 -7302 498504 -7066
rect 497904 -7386 498504 -7302
rect 497904 -7622 498086 -7386
rect 498322 -7622 498504 -7386
rect 497904 -7654 498504 -7622
rect 515904 -6106 516504 13158
rect 522804 705798 523404 705830
rect 522804 705562 522986 705798
rect 523222 705562 523404 705798
rect 522804 705478 523404 705562
rect 522804 705242 522986 705478
rect 523222 705242 523404 705478
rect 522804 668294 523404 705242
rect 522804 668058 522986 668294
rect 523222 668058 523404 668294
rect 522804 632294 523404 668058
rect 522804 632058 522986 632294
rect 523222 632058 523404 632294
rect 522804 596294 523404 632058
rect 522804 596058 522986 596294
rect 523222 596058 523404 596294
rect 522804 560294 523404 596058
rect 522804 560058 522986 560294
rect 523222 560058 523404 560294
rect 522804 524294 523404 560058
rect 522804 524058 522986 524294
rect 523222 524058 523404 524294
rect 522804 488294 523404 524058
rect 522804 488058 522986 488294
rect 523222 488058 523404 488294
rect 522804 452294 523404 488058
rect 522804 452058 522986 452294
rect 523222 452058 523404 452294
rect 522804 416294 523404 452058
rect 522804 416058 522986 416294
rect 523222 416058 523404 416294
rect 522804 380294 523404 416058
rect 522804 380058 522986 380294
rect 523222 380058 523404 380294
rect 522804 344294 523404 380058
rect 522804 344058 522986 344294
rect 523222 344058 523404 344294
rect 522804 308294 523404 344058
rect 522804 308058 522986 308294
rect 523222 308058 523404 308294
rect 522804 272294 523404 308058
rect 522804 272058 522986 272294
rect 523222 272058 523404 272294
rect 522804 236294 523404 272058
rect 522804 236058 522986 236294
rect 523222 236058 523404 236294
rect 522804 200294 523404 236058
rect 522804 200058 522986 200294
rect 523222 200058 523404 200294
rect 522804 164294 523404 200058
rect 522804 164058 522986 164294
rect 523222 164058 523404 164294
rect 522804 128294 523404 164058
rect 522804 128058 522986 128294
rect 523222 128058 523404 128294
rect 522804 92294 523404 128058
rect 522804 92058 522986 92294
rect 523222 92058 523404 92294
rect 522804 56294 523404 92058
rect 522804 56058 522986 56294
rect 523222 56058 523404 56294
rect 522804 20294 523404 56058
rect 522804 20058 522986 20294
rect 523222 20058 523404 20294
rect 522804 -1306 523404 20058
rect 522804 -1542 522986 -1306
rect 523222 -1542 523404 -1306
rect 522804 -1626 523404 -1542
rect 522804 -1862 522986 -1626
rect 523222 -1862 523404 -1626
rect 522804 -1894 523404 -1862
rect 526504 671994 527104 707162
rect 526504 671758 526686 671994
rect 526922 671758 527104 671994
rect 526504 635994 527104 671758
rect 526504 635758 526686 635994
rect 526922 635758 527104 635994
rect 526504 599994 527104 635758
rect 526504 599758 526686 599994
rect 526922 599758 527104 599994
rect 526504 563994 527104 599758
rect 526504 563758 526686 563994
rect 526922 563758 527104 563994
rect 526504 527994 527104 563758
rect 526504 527758 526686 527994
rect 526922 527758 527104 527994
rect 526504 491994 527104 527758
rect 526504 491758 526686 491994
rect 526922 491758 527104 491994
rect 526504 455994 527104 491758
rect 526504 455758 526686 455994
rect 526922 455758 527104 455994
rect 526504 419994 527104 455758
rect 526504 419758 526686 419994
rect 526922 419758 527104 419994
rect 526504 383994 527104 419758
rect 526504 383758 526686 383994
rect 526922 383758 527104 383994
rect 526504 347994 527104 383758
rect 526504 347758 526686 347994
rect 526922 347758 527104 347994
rect 526504 311994 527104 347758
rect 526504 311758 526686 311994
rect 526922 311758 527104 311994
rect 526504 275994 527104 311758
rect 526504 275758 526686 275994
rect 526922 275758 527104 275994
rect 526504 239994 527104 275758
rect 526504 239758 526686 239994
rect 526922 239758 527104 239994
rect 526504 203994 527104 239758
rect 526504 203758 526686 203994
rect 526922 203758 527104 203994
rect 526504 167994 527104 203758
rect 526504 167758 526686 167994
rect 526922 167758 527104 167994
rect 526504 131994 527104 167758
rect 526504 131758 526686 131994
rect 526922 131758 527104 131994
rect 526504 95994 527104 131758
rect 526504 95758 526686 95994
rect 526922 95758 527104 95994
rect 526504 59994 527104 95758
rect 526504 59758 526686 59994
rect 526922 59758 527104 59994
rect 526504 23994 527104 59758
rect 526504 23758 526686 23994
rect 526922 23758 527104 23994
rect 526504 -3226 527104 23758
rect 526504 -3462 526686 -3226
rect 526922 -3462 527104 -3226
rect 526504 -3546 527104 -3462
rect 526504 -3782 526686 -3546
rect 526922 -3782 527104 -3546
rect 526504 -3814 527104 -3782
rect 530204 675694 530804 709082
rect 530204 675458 530386 675694
rect 530622 675458 530804 675694
rect 530204 639694 530804 675458
rect 530204 639458 530386 639694
rect 530622 639458 530804 639694
rect 530204 603694 530804 639458
rect 530204 603458 530386 603694
rect 530622 603458 530804 603694
rect 530204 567694 530804 603458
rect 530204 567458 530386 567694
rect 530622 567458 530804 567694
rect 530204 531694 530804 567458
rect 530204 531458 530386 531694
rect 530622 531458 530804 531694
rect 530204 495694 530804 531458
rect 530204 495458 530386 495694
rect 530622 495458 530804 495694
rect 530204 459694 530804 495458
rect 530204 459458 530386 459694
rect 530622 459458 530804 459694
rect 530204 423694 530804 459458
rect 530204 423458 530386 423694
rect 530622 423458 530804 423694
rect 530204 387694 530804 423458
rect 530204 387458 530386 387694
rect 530622 387458 530804 387694
rect 530204 351694 530804 387458
rect 530204 351458 530386 351694
rect 530622 351458 530804 351694
rect 530204 315694 530804 351458
rect 530204 315458 530386 315694
rect 530622 315458 530804 315694
rect 530204 279694 530804 315458
rect 530204 279458 530386 279694
rect 530622 279458 530804 279694
rect 530204 243694 530804 279458
rect 530204 243458 530386 243694
rect 530622 243458 530804 243694
rect 530204 207694 530804 243458
rect 530204 207458 530386 207694
rect 530622 207458 530804 207694
rect 530204 171694 530804 207458
rect 530204 171458 530386 171694
rect 530622 171458 530804 171694
rect 530204 135694 530804 171458
rect 530204 135458 530386 135694
rect 530622 135458 530804 135694
rect 530204 99694 530804 135458
rect 530204 99458 530386 99694
rect 530622 99458 530804 99694
rect 530204 63694 530804 99458
rect 530204 63458 530386 63694
rect 530622 63458 530804 63694
rect 530204 27694 530804 63458
rect 530204 27458 530386 27694
rect 530622 27458 530804 27694
rect 530204 -5146 530804 27458
rect 530204 -5382 530386 -5146
rect 530622 -5382 530804 -5146
rect 530204 -5466 530804 -5382
rect 530204 -5702 530386 -5466
rect 530622 -5702 530804 -5466
rect 530204 -5734 530804 -5702
rect 533904 679394 534504 711002
rect 551904 710598 552504 711590
rect 551904 710362 552086 710598
rect 552322 710362 552504 710598
rect 551904 710278 552504 710362
rect 551904 710042 552086 710278
rect 552322 710042 552504 710278
rect 548204 708678 548804 709670
rect 548204 708442 548386 708678
rect 548622 708442 548804 708678
rect 548204 708358 548804 708442
rect 548204 708122 548386 708358
rect 548622 708122 548804 708358
rect 544504 706758 545104 707750
rect 544504 706522 544686 706758
rect 544922 706522 545104 706758
rect 544504 706438 545104 706522
rect 544504 706202 544686 706438
rect 544922 706202 545104 706438
rect 533904 679158 534086 679394
rect 534322 679158 534504 679394
rect 533904 643394 534504 679158
rect 533904 643158 534086 643394
rect 534322 643158 534504 643394
rect 533904 607394 534504 643158
rect 533904 607158 534086 607394
rect 534322 607158 534504 607394
rect 533904 571394 534504 607158
rect 533904 571158 534086 571394
rect 534322 571158 534504 571394
rect 533904 535394 534504 571158
rect 533904 535158 534086 535394
rect 534322 535158 534504 535394
rect 533904 499394 534504 535158
rect 533904 499158 534086 499394
rect 534322 499158 534504 499394
rect 533904 463394 534504 499158
rect 533904 463158 534086 463394
rect 534322 463158 534504 463394
rect 533904 427394 534504 463158
rect 533904 427158 534086 427394
rect 534322 427158 534504 427394
rect 533904 391394 534504 427158
rect 533904 391158 534086 391394
rect 534322 391158 534504 391394
rect 533904 355394 534504 391158
rect 533904 355158 534086 355394
rect 534322 355158 534504 355394
rect 533904 319394 534504 355158
rect 533904 319158 534086 319394
rect 534322 319158 534504 319394
rect 533904 283394 534504 319158
rect 533904 283158 534086 283394
rect 534322 283158 534504 283394
rect 533904 247394 534504 283158
rect 533904 247158 534086 247394
rect 534322 247158 534504 247394
rect 533904 211394 534504 247158
rect 533904 211158 534086 211394
rect 534322 211158 534504 211394
rect 533904 175394 534504 211158
rect 533904 175158 534086 175394
rect 534322 175158 534504 175394
rect 533904 139394 534504 175158
rect 533904 139158 534086 139394
rect 534322 139158 534504 139394
rect 533904 103394 534504 139158
rect 533904 103158 534086 103394
rect 534322 103158 534504 103394
rect 533904 67394 534504 103158
rect 533904 67158 534086 67394
rect 534322 67158 534504 67394
rect 533904 31394 534504 67158
rect 533904 31158 534086 31394
rect 534322 31158 534504 31394
rect 515904 -6342 516086 -6106
rect 516322 -6342 516504 -6106
rect 515904 -6426 516504 -6342
rect 515904 -6662 516086 -6426
rect 516322 -6662 516504 -6426
rect 515904 -7654 516504 -6662
rect 533904 -7066 534504 31158
rect 540804 704838 541404 705830
rect 540804 704602 540986 704838
rect 541222 704602 541404 704838
rect 540804 704518 541404 704602
rect 540804 704282 540986 704518
rect 541222 704282 541404 704518
rect 540804 686294 541404 704282
rect 540804 686058 540986 686294
rect 541222 686058 541404 686294
rect 540804 650294 541404 686058
rect 540804 650058 540986 650294
rect 541222 650058 541404 650294
rect 540804 614294 541404 650058
rect 540804 614058 540986 614294
rect 541222 614058 541404 614294
rect 540804 578294 541404 614058
rect 540804 578058 540986 578294
rect 541222 578058 541404 578294
rect 540804 542294 541404 578058
rect 540804 542058 540986 542294
rect 541222 542058 541404 542294
rect 540804 506294 541404 542058
rect 540804 506058 540986 506294
rect 541222 506058 541404 506294
rect 540804 470294 541404 506058
rect 540804 470058 540986 470294
rect 541222 470058 541404 470294
rect 540804 434294 541404 470058
rect 540804 434058 540986 434294
rect 541222 434058 541404 434294
rect 540804 398294 541404 434058
rect 540804 398058 540986 398294
rect 541222 398058 541404 398294
rect 540804 362294 541404 398058
rect 540804 362058 540986 362294
rect 541222 362058 541404 362294
rect 540804 326294 541404 362058
rect 540804 326058 540986 326294
rect 541222 326058 541404 326294
rect 540804 290294 541404 326058
rect 540804 290058 540986 290294
rect 541222 290058 541404 290294
rect 540804 254294 541404 290058
rect 540804 254058 540986 254294
rect 541222 254058 541404 254294
rect 540804 218294 541404 254058
rect 540804 218058 540986 218294
rect 541222 218058 541404 218294
rect 540804 182294 541404 218058
rect 540804 182058 540986 182294
rect 541222 182058 541404 182294
rect 540804 146294 541404 182058
rect 540804 146058 540986 146294
rect 541222 146058 541404 146294
rect 540804 110294 541404 146058
rect 540804 110058 540986 110294
rect 541222 110058 541404 110294
rect 540804 74294 541404 110058
rect 540804 74058 540986 74294
rect 541222 74058 541404 74294
rect 540804 38294 541404 74058
rect 540804 38058 540986 38294
rect 541222 38058 541404 38294
rect 540804 2294 541404 38058
rect 540804 2058 540986 2294
rect 541222 2058 541404 2294
rect 540804 -346 541404 2058
rect 540804 -582 540986 -346
rect 541222 -582 541404 -346
rect 540804 -666 541404 -582
rect 540804 -902 540986 -666
rect 541222 -902 541404 -666
rect 540804 -1894 541404 -902
rect 544504 689994 545104 706202
rect 544504 689758 544686 689994
rect 544922 689758 545104 689994
rect 544504 653994 545104 689758
rect 544504 653758 544686 653994
rect 544922 653758 545104 653994
rect 544504 617994 545104 653758
rect 544504 617758 544686 617994
rect 544922 617758 545104 617994
rect 544504 581994 545104 617758
rect 544504 581758 544686 581994
rect 544922 581758 545104 581994
rect 544504 545994 545104 581758
rect 544504 545758 544686 545994
rect 544922 545758 545104 545994
rect 544504 509994 545104 545758
rect 544504 509758 544686 509994
rect 544922 509758 545104 509994
rect 544504 473994 545104 509758
rect 544504 473758 544686 473994
rect 544922 473758 545104 473994
rect 544504 437994 545104 473758
rect 544504 437758 544686 437994
rect 544922 437758 545104 437994
rect 544504 401994 545104 437758
rect 544504 401758 544686 401994
rect 544922 401758 545104 401994
rect 544504 365994 545104 401758
rect 544504 365758 544686 365994
rect 544922 365758 545104 365994
rect 544504 329994 545104 365758
rect 544504 329758 544686 329994
rect 544922 329758 545104 329994
rect 544504 293994 545104 329758
rect 544504 293758 544686 293994
rect 544922 293758 545104 293994
rect 544504 257994 545104 293758
rect 544504 257758 544686 257994
rect 544922 257758 545104 257994
rect 544504 221994 545104 257758
rect 544504 221758 544686 221994
rect 544922 221758 545104 221994
rect 544504 185994 545104 221758
rect 544504 185758 544686 185994
rect 544922 185758 545104 185994
rect 544504 149994 545104 185758
rect 544504 149758 544686 149994
rect 544922 149758 545104 149994
rect 544504 113994 545104 149758
rect 544504 113758 544686 113994
rect 544922 113758 545104 113994
rect 544504 77994 545104 113758
rect 544504 77758 544686 77994
rect 544922 77758 545104 77994
rect 544504 41994 545104 77758
rect 544504 41758 544686 41994
rect 544922 41758 545104 41994
rect 544504 5994 545104 41758
rect 544504 5758 544686 5994
rect 544922 5758 545104 5994
rect 544504 -2266 545104 5758
rect 544504 -2502 544686 -2266
rect 544922 -2502 545104 -2266
rect 544504 -2586 545104 -2502
rect 544504 -2822 544686 -2586
rect 544922 -2822 545104 -2586
rect 544504 -3814 545104 -2822
rect 548204 693694 548804 708122
rect 548204 693458 548386 693694
rect 548622 693458 548804 693694
rect 548204 657694 548804 693458
rect 548204 657458 548386 657694
rect 548622 657458 548804 657694
rect 548204 621694 548804 657458
rect 548204 621458 548386 621694
rect 548622 621458 548804 621694
rect 548204 585694 548804 621458
rect 548204 585458 548386 585694
rect 548622 585458 548804 585694
rect 548204 549694 548804 585458
rect 548204 549458 548386 549694
rect 548622 549458 548804 549694
rect 548204 513694 548804 549458
rect 548204 513458 548386 513694
rect 548622 513458 548804 513694
rect 548204 477694 548804 513458
rect 548204 477458 548386 477694
rect 548622 477458 548804 477694
rect 548204 441694 548804 477458
rect 548204 441458 548386 441694
rect 548622 441458 548804 441694
rect 548204 405694 548804 441458
rect 548204 405458 548386 405694
rect 548622 405458 548804 405694
rect 548204 369694 548804 405458
rect 548204 369458 548386 369694
rect 548622 369458 548804 369694
rect 548204 333694 548804 369458
rect 548204 333458 548386 333694
rect 548622 333458 548804 333694
rect 548204 297694 548804 333458
rect 548204 297458 548386 297694
rect 548622 297458 548804 297694
rect 548204 261694 548804 297458
rect 548204 261458 548386 261694
rect 548622 261458 548804 261694
rect 548204 225694 548804 261458
rect 548204 225458 548386 225694
rect 548622 225458 548804 225694
rect 548204 189694 548804 225458
rect 548204 189458 548386 189694
rect 548622 189458 548804 189694
rect 548204 153694 548804 189458
rect 548204 153458 548386 153694
rect 548622 153458 548804 153694
rect 548204 117694 548804 153458
rect 548204 117458 548386 117694
rect 548622 117458 548804 117694
rect 548204 81694 548804 117458
rect 548204 81458 548386 81694
rect 548622 81458 548804 81694
rect 548204 45694 548804 81458
rect 548204 45458 548386 45694
rect 548622 45458 548804 45694
rect 548204 9694 548804 45458
rect 548204 9458 548386 9694
rect 548622 9458 548804 9694
rect 548204 -4186 548804 9458
rect 548204 -4422 548386 -4186
rect 548622 -4422 548804 -4186
rect 548204 -4506 548804 -4422
rect 548204 -4742 548386 -4506
rect 548622 -4742 548804 -4506
rect 548204 -5734 548804 -4742
rect 551904 697394 552504 710042
rect 569904 711558 570504 711590
rect 569904 711322 570086 711558
rect 570322 711322 570504 711558
rect 569904 711238 570504 711322
rect 569904 711002 570086 711238
rect 570322 711002 570504 711238
rect 566204 709638 566804 709670
rect 566204 709402 566386 709638
rect 566622 709402 566804 709638
rect 566204 709318 566804 709402
rect 566204 709082 566386 709318
rect 566622 709082 566804 709318
rect 562504 707718 563104 707750
rect 562504 707482 562686 707718
rect 562922 707482 563104 707718
rect 562504 707398 563104 707482
rect 562504 707162 562686 707398
rect 562922 707162 563104 707398
rect 551904 697158 552086 697394
rect 552322 697158 552504 697394
rect 551904 661394 552504 697158
rect 551904 661158 552086 661394
rect 552322 661158 552504 661394
rect 551904 625394 552504 661158
rect 551904 625158 552086 625394
rect 552322 625158 552504 625394
rect 551904 589394 552504 625158
rect 551904 589158 552086 589394
rect 552322 589158 552504 589394
rect 551904 553394 552504 589158
rect 551904 553158 552086 553394
rect 552322 553158 552504 553394
rect 551904 517394 552504 553158
rect 551904 517158 552086 517394
rect 552322 517158 552504 517394
rect 551904 481394 552504 517158
rect 551904 481158 552086 481394
rect 552322 481158 552504 481394
rect 551904 445394 552504 481158
rect 551904 445158 552086 445394
rect 552322 445158 552504 445394
rect 551904 409394 552504 445158
rect 551904 409158 552086 409394
rect 552322 409158 552504 409394
rect 551904 373394 552504 409158
rect 551904 373158 552086 373394
rect 552322 373158 552504 373394
rect 551904 337394 552504 373158
rect 551904 337158 552086 337394
rect 552322 337158 552504 337394
rect 551904 301394 552504 337158
rect 551904 301158 552086 301394
rect 552322 301158 552504 301394
rect 551904 265394 552504 301158
rect 551904 265158 552086 265394
rect 552322 265158 552504 265394
rect 551904 229394 552504 265158
rect 551904 229158 552086 229394
rect 552322 229158 552504 229394
rect 551904 193394 552504 229158
rect 551904 193158 552086 193394
rect 552322 193158 552504 193394
rect 551904 157394 552504 193158
rect 551904 157158 552086 157394
rect 552322 157158 552504 157394
rect 551904 121394 552504 157158
rect 551904 121158 552086 121394
rect 552322 121158 552504 121394
rect 551904 85394 552504 121158
rect 551904 85158 552086 85394
rect 552322 85158 552504 85394
rect 551904 49394 552504 85158
rect 551904 49158 552086 49394
rect 552322 49158 552504 49394
rect 551904 13394 552504 49158
rect 551904 13158 552086 13394
rect 552322 13158 552504 13394
rect 533904 -7302 534086 -7066
rect 534322 -7302 534504 -7066
rect 533904 -7386 534504 -7302
rect 533904 -7622 534086 -7386
rect 534322 -7622 534504 -7386
rect 533904 -7654 534504 -7622
rect 551904 -6106 552504 13158
rect 558804 705798 559404 705830
rect 558804 705562 558986 705798
rect 559222 705562 559404 705798
rect 558804 705478 559404 705562
rect 558804 705242 558986 705478
rect 559222 705242 559404 705478
rect 558804 668294 559404 705242
rect 558804 668058 558986 668294
rect 559222 668058 559404 668294
rect 558804 632294 559404 668058
rect 558804 632058 558986 632294
rect 559222 632058 559404 632294
rect 558804 596294 559404 632058
rect 558804 596058 558986 596294
rect 559222 596058 559404 596294
rect 558804 560294 559404 596058
rect 558804 560058 558986 560294
rect 559222 560058 559404 560294
rect 558804 524294 559404 560058
rect 558804 524058 558986 524294
rect 559222 524058 559404 524294
rect 558804 488294 559404 524058
rect 558804 488058 558986 488294
rect 559222 488058 559404 488294
rect 558804 452294 559404 488058
rect 558804 452058 558986 452294
rect 559222 452058 559404 452294
rect 558804 416294 559404 452058
rect 558804 416058 558986 416294
rect 559222 416058 559404 416294
rect 558804 380294 559404 416058
rect 558804 380058 558986 380294
rect 559222 380058 559404 380294
rect 558804 344294 559404 380058
rect 558804 344058 558986 344294
rect 559222 344058 559404 344294
rect 558804 308294 559404 344058
rect 558804 308058 558986 308294
rect 559222 308058 559404 308294
rect 558804 272294 559404 308058
rect 558804 272058 558986 272294
rect 559222 272058 559404 272294
rect 558804 236294 559404 272058
rect 558804 236058 558986 236294
rect 559222 236058 559404 236294
rect 558804 200294 559404 236058
rect 558804 200058 558986 200294
rect 559222 200058 559404 200294
rect 558804 164294 559404 200058
rect 558804 164058 558986 164294
rect 559222 164058 559404 164294
rect 558804 128294 559404 164058
rect 558804 128058 558986 128294
rect 559222 128058 559404 128294
rect 558804 92294 559404 128058
rect 558804 92058 558986 92294
rect 559222 92058 559404 92294
rect 558804 56294 559404 92058
rect 558804 56058 558986 56294
rect 559222 56058 559404 56294
rect 558804 20294 559404 56058
rect 558804 20058 558986 20294
rect 559222 20058 559404 20294
rect 558804 -1306 559404 20058
rect 558804 -1542 558986 -1306
rect 559222 -1542 559404 -1306
rect 558804 -1626 559404 -1542
rect 558804 -1862 558986 -1626
rect 559222 -1862 559404 -1626
rect 558804 -1894 559404 -1862
rect 562504 671994 563104 707162
rect 562504 671758 562686 671994
rect 562922 671758 563104 671994
rect 562504 635994 563104 671758
rect 562504 635758 562686 635994
rect 562922 635758 563104 635994
rect 562504 599994 563104 635758
rect 562504 599758 562686 599994
rect 562922 599758 563104 599994
rect 562504 563994 563104 599758
rect 562504 563758 562686 563994
rect 562922 563758 563104 563994
rect 562504 527994 563104 563758
rect 562504 527758 562686 527994
rect 562922 527758 563104 527994
rect 562504 491994 563104 527758
rect 562504 491758 562686 491994
rect 562922 491758 563104 491994
rect 562504 455994 563104 491758
rect 562504 455758 562686 455994
rect 562922 455758 563104 455994
rect 562504 419994 563104 455758
rect 562504 419758 562686 419994
rect 562922 419758 563104 419994
rect 562504 383994 563104 419758
rect 562504 383758 562686 383994
rect 562922 383758 563104 383994
rect 562504 347994 563104 383758
rect 562504 347758 562686 347994
rect 562922 347758 563104 347994
rect 562504 311994 563104 347758
rect 562504 311758 562686 311994
rect 562922 311758 563104 311994
rect 562504 275994 563104 311758
rect 562504 275758 562686 275994
rect 562922 275758 563104 275994
rect 562504 239994 563104 275758
rect 562504 239758 562686 239994
rect 562922 239758 563104 239994
rect 562504 203994 563104 239758
rect 562504 203758 562686 203994
rect 562922 203758 563104 203994
rect 562504 167994 563104 203758
rect 562504 167758 562686 167994
rect 562922 167758 563104 167994
rect 562504 131994 563104 167758
rect 562504 131758 562686 131994
rect 562922 131758 563104 131994
rect 562504 95994 563104 131758
rect 562504 95758 562686 95994
rect 562922 95758 563104 95994
rect 562504 59994 563104 95758
rect 562504 59758 562686 59994
rect 562922 59758 563104 59994
rect 562504 23994 563104 59758
rect 562504 23758 562686 23994
rect 562922 23758 563104 23994
rect 562504 -3226 563104 23758
rect 562504 -3462 562686 -3226
rect 562922 -3462 563104 -3226
rect 562504 -3546 563104 -3462
rect 562504 -3782 562686 -3546
rect 562922 -3782 563104 -3546
rect 562504 -3814 563104 -3782
rect 566204 675694 566804 709082
rect 566204 675458 566386 675694
rect 566622 675458 566804 675694
rect 566204 639694 566804 675458
rect 566204 639458 566386 639694
rect 566622 639458 566804 639694
rect 566204 603694 566804 639458
rect 566204 603458 566386 603694
rect 566622 603458 566804 603694
rect 566204 567694 566804 603458
rect 566204 567458 566386 567694
rect 566622 567458 566804 567694
rect 566204 531694 566804 567458
rect 566204 531458 566386 531694
rect 566622 531458 566804 531694
rect 566204 495694 566804 531458
rect 566204 495458 566386 495694
rect 566622 495458 566804 495694
rect 566204 459694 566804 495458
rect 566204 459458 566386 459694
rect 566622 459458 566804 459694
rect 566204 423694 566804 459458
rect 566204 423458 566386 423694
rect 566622 423458 566804 423694
rect 566204 387694 566804 423458
rect 566204 387458 566386 387694
rect 566622 387458 566804 387694
rect 566204 351694 566804 387458
rect 566204 351458 566386 351694
rect 566622 351458 566804 351694
rect 566204 315694 566804 351458
rect 566204 315458 566386 315694
rect 566622 315458 566804 315694
rect 566204 279694 566804 315458
rect 566204 279458 566386 279694
rect 566622 279458 566804 279694
rect 566204 243694 566804 279458
rect 566204 243458 566386 243694
rect 566622 243458 566804 243694
rect 566204 207694 566804 243458
rect 566204 207458 566386 207694
rect 566622 207458 566804 207694
rect 566204 171694 566804 207458
rect 566204 171458 566386 171694
rect 566622 171458 566804 171694
rect 566204 135694 566804 171458
rect 566204 135458 566386 135694
rect 566622 135458 566804 135694
rect 566204 99694 566804 135458
rect 566204 99458 566386 99694
rect 566622 99458 566804 99694
rect 566204 63694 566804 99458
rect 566204 63458 566386 63694
rect 566622 63458 566804 63694
rect 566204 27694 566804 63458
rect 566204 27458 566386 27694
rect 566622 27458 566804 27694
rect 566204 -5146 566804 27458
rect 566204 -5382 566386 -5146
rect 566622 -5382 566804 -5146
rect 566204 -5466 566804 -5382
rect 566204 -5702 566386 -5466
rect 566622 -5702 566804 -5466
rect 566204 -5734 566804 -5702
rect 569904 679394 570504 711002
rect 592030 711558 592650 711590
rect 592030 711322 592062 711558
rect 592298 711322 592382 711558
rect 592618 711322 592650 711558
rect 592030 711238 592650 711322
rect 592030 711002 592062 711238
rect 592298 711002 592382 711238
rect 592618 711002 592650 711238
rect 591070 710598 591690 710630
rect 591070 710362 591102 710598
rect 591338 710362 591422 710598
rect 591658 710362 591690 710598
rect 591070 710278 591690 710362
rect 591070 710042 591102 710278
rect 591338 710042 591422 710278
rect 591658 710042 591690 710278
rect 590110 709638 590730 709670
rect 590110 709402 590142 709638
rect 590378 709402 590462 709638
rect 590698 709402 590730 709638
rect 590110 709318 590730 709402
rect 590110 709082 590142 709318
rect 590378 709082 590462 709318
rect 590698 709082 590730 709318
rect 589150 708678 589770 708710
rect 589150 708442 589182 708678
rect 589418 708442 589502 708678
rect 589738 708442 589770 708678
rect 589150 708358 589770 708442
rect 589150 708122 589182 708358
rect 589418 708122 589502 708358
rect 589738 708122 589770 708358
rect 580504 706758 581104 707750
rect 588190 707718 588810 707750
rect 588190 707482 588222 707718
rect 588458 707482 588542 707718
rect 588778 707482 588810 707718
rect 588190 707398 588810 707482
rect 588190 707162 588222 707398
rect 588458 707162 588542 707398
rect 588778 707162 588810 707398
rect 580504 706522 580686 706758
rect 580922 706522 581104 706758
rect 580504 706438 581104 706522
rect 580504 706202 580686 706438
rect 580922 706202 581104 706438
rect 569904 679158 570086 679394
rect 570322 679158 570504 679394
rect 569904 643394 570504 679158
rect 569904 643158 570086 643394
rect 570322 643158 570504 643394
rect 569904 607394 570504 643158
rect 569904 607158 570086 607394
rect 570322 607158 570504 607394
rect 569904 571394 570504 607158
rect 569904 571158 570086 571394
rect 570322 571158 570504 571394
rect 569904 535394 570504 571158
rect 569904 535158 570086 535394
rect 570322 535158 570504 535394
rect 569904 499394 570504 535158
rect 569904 499158 570086 499394
rect 570322 499158 570504 499394
rect 569904 463394 570504 499158
rect 569904 463158 570086 463394
rect 570322 463158 570504 463394
rect 569904 427394 570504 463158
rect 569904 427158 570086 427394
rect 570322 427158 570504 427394
rect 569904 391394 570504 427158
rect 569904 391158 570086 391394
rect 570322 391158 570504 391394
rect 569904 355394 570504 391158
rect 569904 355158 570086 355394
rect 570322 355158 570504 355394
rect 569904 319394 570504 355158
rect 569904 319158 570086 319394
rect 570322 319158 570504 319394
rect 569904 283394 570504 319158
rect 569904 283158 570086 283394
rect 570322 283158 570504 283394
rect 569904 247394 570504 283158
rect 569904 247158 570086 247394
rect 570322 247158 570504 247394
rect 569904 211394 570504 247158
rect 569904 211158 570086 211394
rect 570322 211158 570504 211394
rect 569904 175394 570504 211158
rect 569904 175158 570086 175394
rect 570322 175158 570504 175394
rect 569904 139394 570504 175158
rect 569904 139158 570086 139394
rect 570322 139158 570504 139394
rect 569904 103394 570504 139158
rect 569904 103158 570086 103394
rect 570322 103158 570504 103394
rect 569904 67394 570504 103158
rect 569904 67158 570086 67394
rect 570322 67158 570504 67394
rect 569904 31394 570504 67158
rect 569904 31158 570086 31394
rect 570322 31158 570504 31394
rect 551904 -6342 552086 -6106
rect 552322 -6342 552504 -6106
rect 551904 -6426 552504 -6342
rect 551904 -6662 552086 -6426
rect 552322 -6662 552504 -6426
rect 551904 -7654 552504 -6662
rect 569904 -7066 570504 31158
rect 576804 704838 577404 705830
rect 576804 704602 576986 704838
rect 577222 704602 577404 704838
rect 576804 704518 577404 704602
rect 576804 704282 576986 704518
rect 577222 704282 577404 704518
rect 576804 686294 577404 704282
rect 576804 686058 576986 686294
rect 577222 686058 577404 686294
rect 576804 650294 577404 686058
rect 576804 650058 576986 650294
rect 577222 650058 577404 650294
rect 576804 614294 577404 650058
rect 576804 614058 576986 614294
rect 577222 614058 577404 614294
rect 576804 578294 577404 614058
rect 576804 578058 576986 578294
rect 577222 578058 577404 578294
rect 576804 542294 577404 578058
rect 576804 542058 576986 542294
rect 577222 542058 577404 542294
rect 576804 506294 577404 542058
rect 576804 506058 576986 506294
rect 577222 506058 577404 506294
rect 576804 470294 577404 506058
rect 576804 470058 576986 470294
rect 577222 470058 577404 470294
rect 576804 434294 577404 470058
rect 576804 434058 576986 434294
rect 577222 434058 577404 434294
rect 576804 398294 577404 434058
rect 576804 398058 576986 398294
rect 577222 398058 577404 398294
rect 576804 362294 577404 398058
rect 576804 362058 576986 362294
rect 577222 362058 577404 362294
rect 576804 326294 577404 362058
rect 576804 326058 576986 326294
rect 577222 326058 577404 326294
rect 576804 290294 577404 326058
rect 576804 290058 576986 290294
rect 577222 290058 577404 290294
rect 576804 254294 577404 290058
rect 576804 254058 576986 254294
rect 577222 254058 577404 254294
rect 576804 218294 577404 254058
rect 576804 218058 576986 218294
rect 577222 218058 577404 218294
rect 576804 182294 577404 218058
rect 576804 182058 576986 182294
rect 577222 182058 577404 182294
rect 576804 146294 577404 182058
rect 576804 146058 576986 146294
rect 577222 146058 577404 146294
rect 576804 110294 577404 146058
rect 576804 110058 576986 110294
rect 577222 110058 577404 110294
rect 576804 74294 577404 110058
rect 576804 74058 576986 74294
rect 577222 74058 577404 74294
rect 576804 38294 577404 74058
rect 576804 38058 576986 38294
rect 577222 38058 577404 38294
rect 576804 2294 577404 38058
rect 576804 2058 576986 2294
rect 577222 2058 577404 2294
rect 576804 -346 577404 2058
rect 576804 -582 576986 -346
rect 577222 -582 577404 -346
rect 576804 -666 577404 -582
rect 576804 -902 576986 -666
rect 577222 -902 577404 -666
rect 576804 -1894 577404 -902
rect 580504 689994 581104 706202
rect 587230 706758 587850 706790
rect 587230 706522 587262 706758
rect 587498 706522 587582 706758
rect 587818 706522 587850 706758
rect 587230 706438 587850 706522
rect 587230 706202 587262 706438
rect 587498 706202 587582 706438
rect 587818 706202 587850 706438
rect 586270 705798 586890 705830
rect 586270 705562 586302 705798
rect 586538 705562 586622 705798
rect 586858 705562 586890 705798
rect 586270 705478 586890 705562
rect 586270 705242 586302 705478
rect 586538 705242 586622 705478
rect 586858 705242 586890 705478
rect 580504 689758 580686 689994
rect 580922 689758 581104 689994
rect 580504 653994 581104 689758
rect 580504 653758 580686 653994
rect 580922 653758 581104 653994
rect 580504 617994 581104 653758
rect 580504 617758 580686 617994
rect 580922 617758 581104 617994
rect 580504 581994 581104 617758
rect 580504 581758 580686 581994
rect 580922 581758 581104 581994
rect 580504 545994 581104 581758
rect 580504 545758 580686 545994
rect 580922 545758 581104 545994
rect 580504 509994 581104 545758
rect 580504 509758 580686 509994
rect 580922 509758 581104 509994
rect 580504 473994 581104 509758
rect 580504 473758 580686 473994
rect 580922 473758 581104 473994
rect 580504 437994 581104 473758
rect 580504 437758 580686 437994
rect 580922 437758 581104 437994
rect 580504 401994 581104 437758
rect 580504 401758 580686 401994
rect 580922 401758 581104 401994
rect 580504 365994 581104 401758
rect 580504 365758 580686 365994
rect 580922 365758 581104 365994
rect 580504 329994 581104 365758
rect 580504 329758 580686 329994
rect 580922 329758 581104 329994
rect 580504 293994 581104 329758
rect 580504 293758 580686 293994
rect 580922 293758 581104 293994
rect 580504 257994 581104 293758
rect 580504 257758 580686 257994
rect 580922 257758 581104 257994
rect 580504 221994 581104 257758
rect 580504 221758 580686 221994
rect 580922 221758 581104 221994
rect 580504 185994 581104 221758
rect 580504 185758 580686 185994
rect 580922 185758 581104 185994
rect 580504 149994 581104 185758
rect 580504 149758 580686 149994
rect 580922 149758 581104 149994
rect 580504 113994 581104 149758
rect 580504 113758 580686 113994
rect 580922 113758 581104 113994
rect 580504 77994 581104 113758
rect 580504 77758 580686 77994
rect 580922 77758 581104 77994
rect 580504 41994 581104 77758
rect 580504 41758 580686 41994
rect 580922 41758 581104 41994
rect 580504 5994 581104 41758
rect 580504 5758 580686 5994
rect 580922 5758 581104 5994
rect 580504 -2266 581104 5758
rect 585310 704838 585930 704870
rect 585310 704602 585342 704838
rect 585578 704602 585662 704838
rect 585898 704602 585930 704838
rect 585310 704518 585930 704602
rect 585310 704282 585342 704518
rect 585578 704282 585662 704518
rect 585898 704282 585930 704518
rect 585310 686294 585930 704282
rect 585310 686058 585342 686294
rect 585578 686058 585662 686294
rect 585898 686058 585930 686294
rect 585310 650294 585930 686058
rect 585310 650058 585342 650294
rect 585578 650058 585662 650294
rect 585898 650058 585930 650294
rect 585310 614294 585930 650058
rect 585310 614058 585342 614294
rect 585578 614058 585662 614294
rect 585898 614058 585930 614294
rect 585310 578294 585930 614058
rect 585310 578058 585342 578294
rect 585578 578058 585662 578294
rect 585898 578058 585930 578294
rect 585310 542294 585930 578058
rect 585310 542058 585342 542294
rect 585578 542058 585662 542294
rect 585898 542058 585930 542294
rect 585310 506294 585930 542058
rect 585310 506058 585342 506294
rect 585578 506058 585662 506294
rect 585898 506058 585930 506294
rect 585310 470294 585930 506058
rect 585310 470058 585342 470294
rect 585578 470058 585662 470294
rect 585898 470058 585930 470294
rect 585310 434294 585930 470058
rect 585310 434058 585342 434294
rect 585578 434058 585662 434294
rect 585898 434058 585930 434294
rect 585310 398294 585930 434058
rect 585310 398058 585342 398294
rect 585578 398058 585662 398294
rect 585898 398058 585930 398294
rect 585310 362294 585930 398058
rect 585310 362058 585342 362294
rect 585578 362058 585662 362294
rect 585898 362058 585930 362294
rect 585310 326294 585930 362058
rect 585310 326058 585342 326294
rect 585578 326058 585662 326294
rect 585898 326058 585930 326294
rect 585310 290294 585930 326058
rect 585310 290058 585342 290294
rect 585578 290058 585662 290294
rect 585898 290058 585930 290294
rect 585310 254294 585930 290058
rect 585310 254058 585342 254294
rect 585578 254058 585662 254294
rect 585898 254058 585930 254294
rect 585310 218294 585930 254058
rect 585310 218058 585342 218294
rect 585578 218058 585662 218294
rect 585898 218058 585930 218294
rect 585310 182294 585930 218058
rect 585310 182058 585342 182294
rect 585578 182058 585662 182294
rect 585898 182058 585930 182294
rect 585310 146294 585930 182058
rect 585310 146058 585342 146294
rect 585578 146058 585662 146294
rect 585898 146058 585930 146294
rect 585310 110294 585930 146058
rect 585310 110058 585342 110294
rect 585578 110058 585662 110294
rect 585898 110058 585930 110294
rect 585310 74294 585930 110058
rect 585310 74058 585342 74294
rect 585578 74058 585662 74294
rect 585898 74058 585930 74294
rect 585310 38294 585930 74058
rect 585310 38058 585342 38294
rect 585578 38058 585662 38294
rect 585898 38058 585930 38294
rect 585310 2294 585930 38058
rect 585310 2058 585342 2294
rect 585578 2058 585662 2294
rect 585898 2058 585930 2294
rect 585310 -346 585930 2058
rect 585310 -582 585342 -346
rect 585578 -582 585662 -346
rect 585898 -582 585930 -346
rect 585310 -666 585930 -582
rect 585310 -902 585342 -666
rect 585578 -902 585662 -666
rect 585898 -902 585930 -666
rect 585310 -934 585930 -902
rect 586270 668294 586890 705242
rect 586270 668058 586302 668294
rect 586538 668058 586622 668294
rect 586858 668058 586890 668294
rect 586270 632294 586890 668058
rect 586270 632058 586302 632294
rect 586538 632058 586622 632294
rect 586858 632058 586890 632294
rect 586270 596294 586890 632058
rect 586270 596058 586302 596294
rect 586538 596058 586622 596294
rect 586858 596058 586890 596294
rect 586270 560294 586890 596058
rect 586270 560058 586302 560294
rect 586538 560058 586622 560294
rect 586858 560058 586890 560294
rect 586270 524294 586890 560058
rect 586270 524058 586302 524294
rect 586538 524058 586622 524294
rect 586858 524058 586890 524294
rect 586270 488294 586890 524058
rect 586270 488058 586302 488294
rect 586538 488058 586622 488294
rect 586858 488058 586890 488294
rect 586270 452294 586890 488058
rect 586270 452058 586302 452294
rect 586538 452058 586622 452294
rect 586858 452058 586890 452294
rect 586270 416294 586890 452058
rect 586270 416058 586302 416294
rect 586538 416058 586622 416294
rect 586858 416058 586890 416294
rect 586270 380294 586890 416058
rect 586270 380058 586302 380294
rect 586538 380058 586622 380294
rect 586858 380058 586890 380294
rect 586270 344294 586890 380058
rect 586270 344058 586302 344294
rect 586538 344058 586622 344294
rect 586858 344058 586890 344294
rect 586270 308294 586890 344058
rect 586270 308058 586302 308294
rect 586538 308058 586622 308294
rect 586858 308058 586890 308294
rect 586270 272294 586890 308058
rect 586270 272058 586302 272294
rect 586538 272058 586622 272294
rect 586858 272058 586890 272294
rect 586270 236294 586890 272058
rect 586270 236058 586302 236294
rect 586538 236058 586622 236294
rect 586858 236058 586890 236294
rect 586270 200294 586890 236058
rect 586270 200058 586302 200294
rect 586538 200058 586622 200294
rect 586858 200058 586890 200294
rect 586270 164294 586890 200058
rect 586270 164058 586302 164294
rect 586538 164058 586622 164294
rect 586858 164058 586890 164294
rect 586270 128294 586890 164058
rect 586270 128058 586302 128294
rect 586538 128058 586622 128294
rect 586858 128058 586890 128294
rect 586270 92294 586890 128058
rect 586270 92058 586302 92294
rect 586538 92058 586622 92294
rect 586858 92058 586890 92294
rect 586270 56294 586890 92058
rect 586270 56058 586302 56294
rect 586538 56058 586622 56294
rect 586858 56058 586890 56294
rect 586270 20294 586890 56058
rect 586270 20058 586302 20294
rect 586538 20058 586622 20294
rect 586858 20058 586890 20294
rect 586270 -1306 586890 20058
rect 586270 -1542 586302 -1306
rect 586538 -1542 586622 -1306
rect 586858 -1542 586890 -1306
rect 586270 -1626 586890 -1542
rect 586270 -1862 586302 -1626
rect 586538 -1862 586622 -1626
rect 586858 -1862 586890 -1626
rect 586270 -1894 586890 -1862
rect 587230 689994 587850 706202
rect 587230 689758 587262 689994
rect 587498 689758 587582 689994
rect 587818 689758 587850 689994
rect 587230 653994 587850 689758
rect 587230 653758 587262 653994
rect 587498 653758 587582 653994
rect 587818 653758 587850 653994
rect 587230 617994 587850 653758
rect 587230 617758 587262 617994
rect 587498 617758 587582 617994
rect 587818 617758 587850 617994
rect 587230 581994 587850 617758
rect 587230 581758 587262 581994
rect 587498 581758 587582 581994
rect 587818 581758 587850 581994
rect 587230 545994 587850 581758
rect 587230 545758 587262 545994
rect 587498 545758 587582 545994
rect 587818 545758 587850 545994
rect 587230 509994 587850 545758
rect 587230 509758 587262 509994
rect 587498 509758 587582 509994
rect 587818 509758 587850 509994
rect 587230 473994 587850 509758
rect 587230 473758 587262 473994
rect 587498 473758 587582 473994
rect 587818 473758 587850 473994
rect 587230 437994 587850 473758
rect 587230 437758 587262 437994
rect 587498 437758 587582 437994
rect 587818 437758 587850 437994
rect 587230 401994 587850 437758
rect 587230 401758 587262 401994
rect 587498 401758 587582 401994
rect 587818 401758 587850 401994
rect 587230 365994 587850 401758
rect 587230 365758 587262 365994
rect 587498 365758 587582 365994
rect 587818 365758 587850 365994
rect 587230 329994 587850 365758
rect 587230 329758 587262 329994
rect 587498 329758 587582 329994
rect 587818 329758 587850 329994
rect 587230 293994 587850 329758
rect 587230 293758 587262 293994
rect 587498 293758 587582 293994
rect 587818 293758 587850 293994
rect 587230 257994 587850 293758
rect 587230 257758 587262 257994
rect 587498 257758 587582 257994
rect 587818 257758 587850 257994
rect 587230 221994 587850 257758
rect 587230 221758 587262 221994
rect 587498 221758 587582 221994
rect 587818 221758 587850 221994
rect 587230 185994 587850 221758
rect 587230 185758 587262 185994
rect 587498 185758 587582 185994
rect 587818 185758 587850 185994
rect 587230 149994 587850 185758
rect 587230 149758 587262 149994
rect 587498 149758 587582 149994
rect 587818 149758 587850 149994
rect 587230 113994 587850 149758
rect 587230 113758 587262 113994
rect 587498 113758 587582 113994
rect 587818 113758 587850 113994
rect 587230 77994 587850 113758
rect 587230 77758 587262 77994
rect 587498 77758 587582 77994
rect 587818 77758 587850 77994
rect 587230 41994 587850 77758
rect 587230 41758 587262 41994
rect 587498 41758 587582 41994
rect 587818 41758 587850 41994
rect 587230 5994 587850 41758
rect 587230 5758 587262 5994
rect 587498 5758 587582 5994
rect 587818 5758 587850 5994
rect 580504 -2502 580686 -2266
rect 580922 -2502 581104 -2266
rect 580504 -2586 581104 -2502
rect 580504 -2822 580686 -2586
rect 580922 -2822 581104 -2586
rect 580504 -3814 581104 -2822
rect 587230 -2266 587850 5758
rect 587230 -2502 587262 -2266
rect 587498 -2502 587582 -2266
rect 587818 -2502 587850 -2266
rect 587230 -2586 587850 -2502
rect 587230 -2822 587262 -2586
rect 587498 -2822 587582 -2586
rect 587818 -2822 587850 -2586
rect 587230 -2854 587850 -2822
rect 588190 671994 588810 707162
rect 588190 671758 588222 671994
rect 588458 671758 588542 671994
rect 588778 671758 588810 671994
rect 588190 635994 588810 671758
rect 588190 635758 588222 635994
rect 588458 635758 588542 635994
rect 588778 635758 588810 635994
rect 588190 599994 588810 635758
rect 588190 599758 588222 599994
rect 588458 599758 588542 599994
rect 588778 599758 588810 599994
rect 588190 563994 588810 599758
rect 588190 563758 588222 563994
rect 588458 563758 588542 563994
rect 588778 563758 588810 563994
rect 588190 527994 588810 563758
rect 588190 527758 588222 527994
rect 588458 527758 588542 527994
rect 588778 527758 588810 527994
rect 588190 491994 588810 527758
rect 588190 491758 588222 491994
rect 588458 491758 588542 491994
rect 588778 491758 588810 491994
rect 588190 455994 588810 491758
rect 588190 455758 588222 455994
rect 588458 455758 588542 455994
rect 588778 455758 588810 455994
rect 588190 419994 588810 455758
rect 588190 419758 588222 419994
rect 588458 419758 588542 419994
rect 588778 419758 588810 419994
rect 588190 383994 588810 419758
rect 588190 383758 588222 383994
rect 588458 383758 588542 383994
rect 588778 383758 588810 383994
rect 588190 347994 588810 383758
rect 588190 347758 588222 347994
rect 588458 347758 588542 347994
rect 588778 347758 588810 347994
rect 588190 311994 588810 347758
rect 588190 311758 588222 311994
rect 588458 311758 588542 311994
rect 588778 311758 588810 311994
rect 588190 275994 588810 311758
rect 588190 275758 588222 275994
rect 588458 275758 588542 275994
rect 588778 275758 588810 275994
rect 588190 239994 588810 275758
rect 588190 239758 588222 239994
rect 588458 239758 588542 239994
rect 588778 239758 588810 239994
rect 588190 203994 588810 239758
rect 588190 203758 588222 203994
rect 588458 203758 588542 203994
rect 588778 203758 588810 203994
rect 588190 167994 588810 203758
rect 588190 167758 588222 167994
rect 588458 167758 588542 167994
rect 588778 167758 588810 167994
rect 588190 131994 588810 167758
rect 588190 131758 588222 131994
rect 588458 131758 588542 131994
rect 588778 131758 588810 131994
rect 588190 95994 588810 131758
rect 588190 95758 588222 95994
rect 588458 95758 588542 95994
rect 588778 95758 588810 95994
rect 588190 59994 588810 95758
rect 588190 59758 588222 59994
rect 588458 59758 588542 59994
rect 588778 59758 588810 59994
rect 588190 23994 588810 59758
rect 588190 23758 588222 23994
rect 588458 23758 588542 23994
rect 588778 23758 588810 23994
rect 588190 -3226 588810 23758
rect 588190 -3462 588222 -3226
rect 588458 -3462 588542 -3226
rect 588778 -3462 588810 -3226
rect 588190 -3546 588810 -3462
rect 588190 -3782 588222 -3546
rect 588458 -3782 588542 -3546
rect 588778 -3782 588810 -3546
rect 588190 -3814 588810 -3782
rect 589150 693694 589770 708122
rect 589150 693458 589182 693694
rect 589418 693458 589502 693694
rect 589738 693458 589770 693694
rect 589150 657694 589770 693458
rect 589150 657458 589182 657694
rect 589418 657458 589502 657694
rect 589738 657458 589770 657694
rect 589150 621694 589770 657458
rect 589150 621458 589182 621694
rect 589418 621458 589502 621694
rect 589738 621458 589770 621694
rect 589150 585694 589770 621458
rect 589150 585458 589182 585694
rect 589418 585458 589502 585694
rect 589738 585458 589770 585694
rect 589150 549694 589770 585458
rect 589150 549458 589182 549694
rect 589418 549458 589502 549694
rect 589738 549458 589770 549694
rect 589150 513694 589770 549458
rect 589150 513458 589182 513694
rect 589418 513458 589502 513694
rect 589738 513458 589770 513694
rect 589150 477694 589770 513458
rect 589150 477458 589182 477694
rect 589418 477458 589502 477694
rect 589738 477458 589770 477694
rect 589150 441694 589770 477458
rect 589150 441458 589182 441694
rect 589418 441458 589502 441694
rect 589738 441458 589770 441694
rect 589150 405694 589770 441458
rect 589150 405458 589182 405694
rect 589418 405458 589502 405694
rect 589738 405458 589770 405694
rect 589150 369694 589770 405458
rect 589150 369458 589182 369694
rect 589418 369458 589502 369694
rect 589738 369458 589770 369694
rect 589150 333694 589770 369458
rect 589150 333458 589182 333694
rect 589418 333458 589502 333694
rect 589738 333458 589770 333694
rect 589150 297694 589770 333458
rect 589150 297458 589182 297694
rect 589418 297458 589502 297694
rect 589738 297458 589770 297694
rect 589150 261694 589770 297458
rect 589150 261458 589182 261694
rect 589418 261458 589502 261694
rect 589738 261458 589770 261694
rect 589150 225694 589770 261458
rect 589150 225458 589182 225694
rect 589418 225458 589502 225694
rect 589738 225458 589770 225694
rect 589150 189694 589770 225458
rect 589150 189458 589182 189694
rect 589418 189458 589502 189694
rect 589738 189458 589770 189694
rect 589150 153694 589770 189458
rect 589150 153458 589182 153694
rect 589418 153458 589502 153694
rect 589738 153458 589770 153694
rect 589150 117694 589770 153458
rect 589150 117458 589182 117694
rect 589418 117458 589502 117694
rect 589738 117458 589770 117694
rect 589150 81694 589770 117458
rect 589150 81458 589182 81694
rect 589418 81458 589502 81694
rect 589738 81458 589770 81694
rect 589150 45694 589770 81458
rect 589150 45458 589182 45694
rect 589418 45458 589502 45694
rect 589738 45458 589770 45694
rect 589150 9694 589770 45458
rect 589150 9458 589182 9694
rect 589418 9458 589502 9694
rect 589738 9458 589770 9694
rect 589150 -4186 589770 9458
rect 589150 -4422 589182 -4186
rect 589418 -4422 589502 -4186
rect 589738 -4422 589770 -4186
rect 589150 -4506 589770 -4422
rect 589150 -4742 589182 -4506
rect 589418 -4742 589502 -4506
rect 589738 -4742 589770 -4506
rect 589150 -4774 589770 -4742
rect 590110 675694 590730 709082
rect 590110 675458 590142 675694
rect 590378 675458 590462 675694
rect 590698 675458 590730 675694
rect 590110 639694 590730 675458
rect 590110 639458 590142 639694
rect 590378 639458 590462 639694
rect 590698 639458 590730 639694
rect 590110 603694 590730 639458
rect 590110 603458 590142 603694
rect 590378 603458 590462 603694
rect 590698 603458 590730 603694
rect 590110 567694 590730 603458
rect 590110 567458 590142 567694
rect 590378 567458 590462 567694
rect 590698 567458 590730 567694
rect 590110 531694 590730 567458
rect 590110 531458 590142 531694
rect 590378 531458 590462 531694
rect 590698 531458 590730 531694
rect 590110 495694 590730 531458
rect 590110 495458 590142 495694
rect 590378 495458 590462 495694
rect 590698 495458 590730 495694
rect 590110 459694 590730 495458
rect 590110 459458 590142 459694
rect 590378 459458 590462 459694
rect 590698 459458 590730 459694
rect 590110 423694 590730 459458
rect 590110 423458 590142 423694
rect 590378 423458 590462 423694
rect 590698 423458 590730 423694
rect 590110 387694 590730 423458
rect 590110 387458 590142 387694
rect 590378 387458 590462 387694
rect 590698 387458 590730 387694
rect 590110 351694 590730 387458
rect 590110 351458 590142 351694
rect 590378 351458 590462 351694
rect 590698 351458 590730 351694
rect 590110 315694 590730 351458
rect 590110 315458 590142 315694
rect 590378 315458 590462 315694
rect 590698 315458 590730 315694
rect 590110 279694 590730 315458
rect 590110 279458 590142 279694
rect 590378 279458 590462 279694
rect 590698 279458 590730 279694
rect 590110 243694 590730 279458
rect 590110 243458 590142 243694
rect 590378 243458 590462 243694
rect 590698 243458 590730 243694
rect 590110 207694 590730 243458
rect 590110 207458 590142 207694
rect 590378 207458 590462 207694
rect 590698 207458 590730 207694
rect 590110 171694 590730 207458
rect 590110 171458 590142 171694
rect 590378 171458 590462 171694
rect 590698 171458 590730 171694
rect 590110 135694 590730 171458
rect 590110 135458 590142 135694
rect 590378 135458 590462 135694
rect 590698 135458 590730 135694
rect 590110 99694 590730 135458
rect 590110 99458 590142 99694
rect 590378 99458 590462 99694
rect 590698 99458 590730 99694
rect 590110 63694 590730 99458
rect 590110 63458 590142 63694
rect 590378 63458 590462 63694
rect 590698 63458 590730 63694
rect 590110 27694 590730 63458
rect 590110 27458 590142 27694
rect 590378 27458 590462 27694
rect 590698 27458 590730 27694
rect 590110 -5146 590730 27458
rect 590110 -5382 590142 -5146
rect 590378 -5382 590462 -5146
rect 590698 -5382 590730 -5146
rect 590110 -5466 590730 -5382
rect 590110 -5702 590142 -5466
rect 590378 -5702 590462 -5466
rect 590698 -5702 590730 -5466
rect 590110 -5734 590730 -5702
rect 591070 697394 591690 710042
rect 591070 697158 591102 697394
rect 591338 697158 591422 697394
rect 591658 697158 591690 697394
rect 591070 661394 591690 697158
rect 591070 661158 591102 661394
rect 591338 661158 591422 661394
rect 591658 661158 591690 661394
rect 591070 625394 591690 661158
rect 591070 625158 591102 625394
rect 591338 625158 591422 625394
rect 591658 625158 591690 625394
rect 591070 589394 591690 625158
rect 591070 589158 591102 589394
rect 591338 589158 591422 589394
rect 591658 589158 591690 589394
rect 591070 553394 591690 589158
rect 591070 553158 591102 553394
rect 591338 553158 591422 553394
rect 591658 553158 591690 553394
rect 591070 517394 591690 553158
rect 591070 517158 591102 517394
rect 591338 517158 591422 517394
rect 591658 517158 591690 517394
rect 591070 481394 591690 517158
rect 591070 481158 591102 481394
rect 591338 481158 591422 481394
rect 591658 481158 591690 481394
rect 591070 445394 591690 481158
rect 591070 445158 591102 445394
rect 591338 445158 591422 445394
rect 591658 445158 591690 445394
rect 591070 409394 591690 445158
rect 591070 409158 591102 409394
rect 591338 409158 591422 409394
rect 591658 409158 591690 409394
rect 591070 373394 591690 409158
rect 591070 373158 591102 373394
rect 591338 373158 591422 373394
rect 591658 373158 591690 373394
rect 591070 337394 591690 373158
rect 591070 337158 591102 337394
rect 591338 337158 591422 337394
rect 591658 337158 591690 337394
rect 591070 301394 591690 337158
rect 591070 301158 591102 301394
rect 591338 301158 591422 301394
rect 591658 301158 591690 301394
rect 591070 265394 591690 301158
rect 591070 265158 591102 265394
rect 591338 265158 591422 265394
rect 591658 265158 591690 265394
rect 591070 229394 591690 265158
rect 591070 229158 591102 229394
rect 591338 229158 591422 229394
rect 591658 229158 591690 229394
rect 591070 193394 591690 229158
rect 591070 193158 591102 193394
rect 591338 193158 591422 193394
rect 591658 193158 591690 193394
rect 591070 157394 591690 193158
rect 591070 157158 591102 157394
rect 591338 157158 591422 157394
rect 591658 157158 591690 157394
rect 591070 121394 591690 157158
rect 591070 121158 591102 121394
rect 591338 121158 591422 121394
rect 591658 121158 591690 121394
rect 591070 85394 591690 121158
rect 591070 85158 591102 85394
rect 591338 85158 591422 85394
rect 591658 85158 591690 85394
rect 591070 49394 591690 85158
rect 591070 49158 591102 49394
rect 591338 49158 591422 49394
rect 591658 49158 591690 49394
rect 591070 13394 591690 49158
rect 591070 13158 591102 13394
rect 591338 13158 591422 13394
rect 591658 13158 591690 13394
rect 591070 -6106 591690 13158
rect 591070 -6342 591102 -6106
rect 591338 -6342 591422 -6106
rect 591658 -6342 591690 -6106
rect 591070 -6426 591690 -6342
rect 591070 -6662 591102 -6426
rect 591338 -6662 591422 -6426
rect 591658 -6662 591690 -6426
rect 591070 -6694 591690 -6662
rect 592030 679394 592650 711002
rect 592030 679158 592062 679394
rect 592298 679158 592382 679394
rect 592618 679158 592650 679394
rect 592030 643394 592650 679158
rect 592030 643158 592062 643394
rect 592298 643158 592382 643394
rect 592618 643158 592650 643394
rect 592030 607394 592650 643158
rect 592030 607158 592062 607394
rect 592298 607158 592382 607394
rect 592618 607158 592650 607394
rect 592030 571394 592650 607158
rect 592030 571158 592062 571394
rect 592298 571158 592382 571394
rect 592618 571158 592650 571394
rect 592030 535394 592650 571158
rect 592030 535158 592062 535394
rect 592298 535158 592382 535394
rect 592618 535158 592650 535394
rect 592030 499394 592650 535158
rect 592030 499158 592062 499394
rect 592298 499158 592382 499394
rect 592618 499158 592650 499394
rect 592030 463394 592650 499158
rect 592030 463158 592062 463394
rect 592298 463158 592382 463394
rect 592618 463158 592650 463394
rect 592030 427394 592650 463158
rect 592030 427158 592062 427394
rect 592298 427158 592382 427394
rect 592618 427158 592650 427394
rect 592030 391394 592650 427158
rect 592030 391158 592062 391394
rect 592298 391158 592382 391394
rect 592618 391158 592650 391394
rect 592030 355394 592650 391158
rect 592030 355158 592062 355394
rect 592298 355158 592382 355394
rect 592618 355158 592650 355394
rect 592030 319394 592650 355158
rect 592030 319158 592062 319394
rect 592298 319158 592382 319394
rect 592618 319158 592650 319394
rect 592030 283394 592650 319158
rect 592030 283158 592062 283394
rect 592298 283158 592382 283394
rect 592618 283158 592650 283394
rect 592030 247394 592650 283158
rect 592030 247158 592062 247394
rect 592298 247158 592382 247394
rect 592618 247158 592650 247394
rect 592030 211394 592650 247158
rect 592030 211158 592062 211394
rect 592298 211158 592382 211394
rect 592618 211158 592650 211394
rect 592030 175394 592650 211158
rect 592030 175158 592062 175394
rect 592298 175158 592382 175394
rect 592618 175158 592650 175394
rect 592030 139394 592650 175158
rect 592030 139158 592062 139394
rect 592298 139158 592382 139394
rect 592618 139158 592650 139394
rect 592030 103394 592650 139158
rect 592030 103158 592062 103394
rect 592298 103158 592382 103394
rect 592618 103158 592650 103394
rect 592030 67394 592650 103158
rect 592030 67158 592062 67394
rect 592298 67158 592382 67394
rect 592618 67158 592650 67394
rect 592030 31394 592650 67158
rect 592030 31158 592062 31394
rect 592298 31158 592382 31394
rect 592618 31158 592650 31394
rect 569904 -7302 570086 -7066
rect 570322 -7302 570504 -7066
rect 569904 -7386 570504 -7302
rect 569904 -7622 570086 -7386
rect 570322 -7622 570504 -7386
rect 569904 -7654 570504 -7622
rect 592030 -7066 592650 31158
rect 592030 -7302 592062 -7066
rect 592298 -7302 592382 -7066
rect 592618 -7302 592650 -7066
rect 592030 -7386 592650 -7302
rect 592030 -7622 592062 -7386
rect 592298 -7622 592382 -7386
rect 592618 -7622 592650 -7386
rect 592030 -7654 592650 -7622
<< via4 >>
rect -8694 711322 -8458 711558
rect -8374 711322 -8138 711558
rect -8694 711002 -8458 711238
rect -8374 711002 -8138 711238
rect -8694 679158 -8458 679394
rect -8374 679158 -8138 679394
rect -8694 643158 -8458 643394
rect -8374 643158 -8138 643394
rect -8694 607158 -8458 607394
rect -8374 607158 -8138 607394
rect -8694 571158 -8458 571394
rect -8374 571158 -8138 571394
rect -8694 535158 -8458 535394
rect -8374 535158 -8138 535394
rect -8694 499158 -8458 499394
rect -8374 499158 -8138 499394
rect -8694 463158 -8458 463394
rect -8374 463158 -8138 463394
rect -8694 427158 -8458 427394
rect -8374 427158 -8138 427394
rect -8694 391158 -8458 391394
rect -8374 391158 -8138 391394
rect -8694 355158 -8458 355394
rect -8374 355158 -8138 355394
rect -8694 319158 -8458 319394
rect -8374 319158 -8138 319394
rect -8694 283158 -8458 283394
rect -8374 283158 -8138 283394
rect -8694 247158 -8458 247394
rect -8374 247158 -8138 247394
rect -8694 211158 -8458 211394
rect -8374 211158 -8138 211394
rect -8694 175158 -8458 175394
rect -8374 175158 -8138 175394
rect -8694 139158 -8458 139394
rect -8374 139158 -8138 139394
rect -8694 103158 -8458 103394
rect -8374 103158 -8138 103394
rect -8694 67158 -8458 67394
rect -8374 67158 -8138 67394
rect -8694 31158 -8458 31394
rect -8374 31158 -8138 31394
rect -7734 710362 -7498 710598
rect -7414 710362 -7178 710598
rect -7734 710042 -7498 710278
rect -7414 710042 -7178 710278
rect 12086 710362 12322 710598
rect 12086 710042 12322 710278
rect -7734 697158 -7498 697394
rect -7414 697158 -7178 697394
rect -7734 661158 -7498 661394
rect -7414 661158 -7178 661394
rect -7734 625158 -7498 625394
rect -7414 625158 -7178 625394
rect -7734 589158 -7498 589394
rect -7414 589158 -7178 589394
rect -7734 553158 -7498 553394
rect -7414 553158 -7178 553394
rect -7734 517158 -7498 517394
rect -7414 517158 -7178 517394
rect -7734 481158 -7498 481394
rect -7414 481158 -7178 481394
rect -7734 445158 -7498 445394
rect -7414 445158 -7178 445394
rect -7734 409158 -7498 409394
rect -7414 409158 -7178 409394
rect -7734 373158 -7498 373394
rect -7414 373158 -7178 373394
rect -7734 337158 -7498 337394
rect -7414 337158 -7178 337394
rect -7734 301158 -7498 301394
rect -7414 301158 -7178 301394
rect -7734 265158 -7498 265394
rect -7414 265158 -7178 265394
rect -7734 229158 -7498 229394
rect -7414 229158 -7178 229394
rect -7734 193158 -7498 193394
rect -7414 193158 -7178 193394
rect -7734 157158 -7498 157394
rect -7414 157158 -7178 157394
rect -7734 121158 -7498 121394
rect -7414 121158 -7178 121394
rect -7734 85158 -7498 85394
rect -7414 85158 -7178 85394
rect -7734 49158 -7498 49394
rect -7414 49158 -7178 49394
rect -7734 13158 -7498 13394
rect -7414 13158 -7178 13394
rect -6774 709402 -6538 709638
rect -6454 709402 -6218 709638
rect -6774 709082 -6538 709318
rect -6454 709082 -6218 709318
rect -6774 675458 -6538 675694
rect -6454 675458 -6218 675694
rect -6774 639458 -6538 639694
rect -6454 639458 -6218 639694
rect -6774 603458 -6538 603694
rect -6454 603458 -6218 603694
rect -6774 567458 -6538 567694
rect -6454 567458 -6218 567694
rect -6774 531458 -6538 531694
rect -6454 531458 -6218 531694
rect -6774 495458 -6538 495694
rect -6454 495458 -6218 495694
rect -6774 459458 -6538 459694
rect -6454 459458 -6218 459694
rect -6774 423458 -6538 423694
rect -6454 423458 -6218 423694
rect -6774 387458 -6538 387694
rect -6454 387458 -6218 387694
rect -6774 351458 -6538 351694
rect -6454 351458 -6218 351694
rect -6774 315458 -6538 315694
rect -6454 315458 -6218 315694
rect -6774 279458 -6538 279694
rect -6454 279458 -6218 279694
rect -6774 243458 -6538 243694
rect -6454 243458 -6218 243694
rect -6774 207458 -6538 207694
rect -6454 207458 -6218 207694
rect -6774 171458 -6538 171694
rect -6454 171458 -6218 171694
rect -6774 135458 -6538 135694
rect -6454 135458 -6218 135694
rect -6774 99458 -6538 99694
rect -6454 99458 -6218 99694
rect -6774 63458 -6538 63694
rect -6454 63458 -6218 63694
rect -6774 27458 -6538 27694
rect -6454 27458 -6218 27694
rect -5814 708442 -5578 708678
rect -5494 708442 -5258 708678
rect -5814 708122 -5578 708358
rect -5494 708122 -5258 708358
rect 8386 708442 8622 708678
rect 8386 708122 8622 708358
rect -5814 693458 -5578 693694
rect -5494 693458 -5258 693694
rect -5814 657458 -5578 657694
rect -5494 657458 -5258 657694
rect -5814 621458 -5578 621694
rect -5494 621458 -5258 621694
rect -5814 585458 -5578 585694
rect -5494 585458 -5258 585694
rect -5814 549458 -5578 549694
rect -5494 549458 -5258 549694
rect -5814 513458 -5578 513694
rect -5494 513458 -5258 513694
rect -5814 477458 -5578 477694
rect -5494 477458 -5258 477694
rect -5814 441458 -5578 441694
rect -5494 441458 -5258 441694
rect -5814 405458 -5578 405694
rect -5494 405458 -5258 405694
rect -5814 369458 -5578 369694
rect -5494 369458 -5258 369694
rect -5814 333458 -5578 333694
rect -5494 333458 -5258 333694
rect -5814 297458 -5578 297694
rect -5494 297458 -5258 297694
rect -5814 261458 -5578 261694
rect -5494 261458 -5258 261694
rect -5814 225458 -5578 225694
rect -5494 225458 -5258 225694
rect -5814 189458 -5578 189694
rect -5494 189458 -5258 189694
rect -5814 153458 -5578 153694
rect -5494 153458 -5258 153694
rect -5814 117458 -5578 117694
rect -5494 117458 -5258 117694
rect -5814 81458 -5578 81694
rect -5494 81458 -5258 81694
rect -5814 45458 -5578 45694
rect -5494 45458 -5258 45694
rect -5814 9458 -5578 9694
rect -5494 9458 -5258 9694
rect -4854 707482 -4618 707718
rect -4534 707482 -4298 707718
rect -4854 707162 -4618 707398
rect -4534 707162 -4298 707398
rect -4854 671758 -4618 671994
rect -4534 671758 -4298 671994
rect -4854 635758 -4618 635994
rect -4534 635758 -4298 635994
rect -4854 599758 -4618 599994
rect -4534 599758 -4298 599994
rect -4854 563758 -4618 563994
rect -4534 563758 -4298 563994
rect -4854 527758 -4618 527994
rect -4534 527758 -4298 527994
rect -4854 491758 -4618 491994
rect -4534 491758 -4298 491994
rect -4854 455758 -4618 455994
rect -4534 455758 -4298 455994
rect -4854 419758 -4618 419994
rect -4534 419758 -4298 419994
rect -4854 383758 -4618 383994
rect -4534 383758 -4298 383994
rect -4854 347758 -4618 347994
rect -4534 347758 -4298 347994
rect -4854 311758 -4618 311994
rect -4534 311758 -4298 311994
rect -4854 275758 -4618 275994
rect -4534 275758 -4298 275994
rect -4854 239758 -4618 239994
rect -4534 239758 -4298 239994
rect -4854 203758 -4618 203994
rect -4534 203758 -4298 203994
rect -4854 167758 -4618 167994
rect -4534 167758 -4298 167994
rect -4854 131758 -4618 131994
rect -4534 131758 -4298 131994
rect -4854 95758 -4618 95994
rect -4534 95758 -4298 95994
rect -4854 59758 -4618 59994
rect -4534 59758 -4298 59994
rect -4854 23758 -4618 23994
rect -4534 23758 -4298 23994
rect -3894 706522 -3658 706758
rect -3574 706522 -3338 706758
rect -3894 706202 -3658 706438
rect -3574 706202 -3338 706438
rect 4686 706522 4922 706758
rect 4686 706202 4922 706438
rect -3894 689758 -3658 689994
rect -3574 689758 -3338 689994
rect -3894 653758 -3658 653994
rect -3574 653758 -3338 653994
rect -3894 617758 -3658 617994
rect -3574 617758 -3338 617994
rect -3894 581758 -3658 581994
rect -3574 581758 -3338 581994
rect -3894 545758 -3658 545994
rect -3574 545758 -3338 545994
rect -3894 509758 -3658 509994
rect -3574 509758 -3338 509994
rect -3894 473758 -3658 473994
rect -3574 473758 -3338 473994
rect -3894 437758 -3658 437994
rect -3574 437758 -3338 437994
rect -3894 401758 -3658 401994
rect -3574 401758 -3338 401994
rect -3894 365758 -3658 365994
rect -3574 365758 -3338 365994
rect -3894 329758 -3658 329994
rect -3574 329758 -3338 329994
rect -3894 293758 -3658 293994
rect -3574 293758 -3338 293994
rect -3894 257758 -3658 257994
rect -3574 257758 -3338 257994
rect -3894 221758 -3658 221994
rect -3574 221758 -3338 221994
rect -3894 185758 -3658 185994
rect -3574 185758 -3338 185994
rect -3894 149758 -3658 149994
rect -3574 149758 -3338 149994
rect -3894 113758 -3658 113994
rect -3574 113758 -3338 113994
rect -3894 77758 -3658 77994
rect -3574 77758 -3338 77994
rect -3894 41758 -3658 41994
rect -3574 41758 -3338 41994
rect -3894 5758 -3658 5994
rect -3574 5758 -3338 5994
rect -2934 705562 -2698 705798
rect -2614 705562 -2378 705798
rect -2934 705242 -2698 705478
rect -2614 705242 -2378 705478
rect -2934 668058 -2698 668294
rect -2614 668058 -2378 668294
rect -2934 632058 -2698 632294
rect -2614 632058 -2378 632294
rect -2934 596058 -2698 596294
rect -2614 596058 -2378 596294
rect -2934 560058 -2698 560294
rect -2614 560058 -2378 560294
rect -2934 524058 -2698 524294
rect -2614 524058 -2378 524294
rect -2934 488058 -2698 488294
rect -2614 488058 -2378 488294
rect -2934 452058 -2698 452294
rect -2614 452058 -2378 452294
rect -2934 416058 -2698 416294
rect -2614 416058 -2378 416294
rect -2934 380058 -2698 380294
rect -2614 380058 -2378 380294
rect -2934 344058 -2698 344294
rect -2614 344058 -2378 344294
rect -2934 308058 -2698 308294
rect -2614 308058 -2378 308294
rect -2934 272058 -2698 272294
rect -2614 272058 -2378 272294
rect -2934 236058 -2698 236294
rect -2614 236058 -2378 236294
rect -2934 200058 -2698 200294
rect -2614 200058 -2378 200294
rect -2934 164058 -2698 164294
rect -2614 164058 -2378 164294
rect -2934 128058 -2698 128294
rect -2614 128058 -2378 128294
rect -2934 92058 -2698 92294
rect -2614 92058 -2378 92294
rect -2934 56058 -2698 56294
rect -2614 56058 -2378 56294
rect -2934 20058 -2698 20294
rect -2614 20058 -2378 20294
rect -1974 704602 -1738 704838
rect -1654 704602 -1418 704838
rect -1974 704282 -1738 704518
rect -1654 704282 -1418 704518
rect -1974 686058 -1738 686294
rect -1654 686058 -1418 686294
rect -1974 650058 -1738 650294
rect -1654 650058 -1418 650294
rect -1974 614058 -1738 614294
rect -1654 614058 -1418 614294
rect -1974 578058 -1738 578294
rect -1654 578058 -1418 578294
rect -1974 542058 -1738 542294
rect -1654 542058 -1418 542294
rect -1974 506058 -1738 506294
rect -1654 506058 -1418 506294
rect -1974 470058 -1738 470294
rect -1654 470058 -1418 470294
rect -1974 434058 -1738 434294
rect -1654 434058 -1418 434294
rect -1974 398058 -1738 398294
rect -1654 398058 -1418 398294
rect -1974 362058 -1738 362294
rect -1654 362058 -1418 362294
rect -1974 326058 -1738 326294
rect -1654 326058 -1418 326294
rect -1974 290058 -1738 290294
rect -1654 290058 -1418 290294
rect -1974 254058 -1738 254294
rect -1654 254058 -1418 254294
rect -1974 218058 -1738 218294
rect -1654 218058 -1418 218294
rect -1974 182058 -1738 182294
rect -1654 182058 -1418 182294
rect -1974 146058 -1738 146294
rect -1654 146058 -1418 146294
rect -1974 110058 -1738 110294
rect -1654 110058 -1418 110294
rect -1974 74058 -1738 74294
rect -1654 74058 -1418 74294
rect -1974 38058 -1738 38294
rect -1654 38058 -1418 38294
rect -1974 2058 -1738 2294
rect -1654 2058 -1418 2294
rect -1974 -582 -1738 -346
rect -1654 -582 -1418 -346
rect -1974 -902 -1738 -666
rect -1654 -902 -1418 -666
rect 986 704602 1222 704838
rect 986 704282 1222 704518
rect 986 686058 1222 686294
rect 986 650058 1222 650294
rect 986 614058 1222 614294
rect 986 578058 1222 578294
rect 986 542058 1222 542294
rect 986 506058 1222 506294
rect 986 470058 1222 470294
rect 986 434058 1222 434294
rect 986 398058 1222 398294
rect 986 362058 1222 362294
rect 986 326058 1222 326294
rect 986 290058 1222 290294
rect 986 254058 1222 254294
rect 986 218058 1222 218294
rect 986 182058 1222 182294
rect 986 146058 1222 146294
rect 986 110058 1222 110294
rect 986 74058 1222 74294
rect 986 38058 1222 38294
rect 986 2058 1222 2294
rect 986 -582 1222 -346
rect 986 -902 1222 -666
rect -2934 -1542 -2698 -1306
rect -2614 -1542 -2378 -1306
rect -2934 -1862 -2698 -1626
rect -2614 -1862 -2378 -1626
rect 4686 689758 4922 689994
rect 4686 653758 4922 653994
rect 4686 617758 4922 617994
rect 4686 581758 4922 581994
rect 4686 545758 4922 545994
rect 4686 509758 4922 509994
rect 4686 473758 4922 473994
rect 4686 437758 4922 437994
rect 4686 401758 4922 401994
rect 4686 365758 4922 365994
rect 4686 329758 4922 329994
rect 4686 293758 4922 293994
rect 4686 257758 4922 257994
rect 4686 221758 4922 221994
rect 4686 185758 4922 185994
rect 4686 149758 4922 149994
rect 4686 113758 4922 113994
rect 4686 77758 4922 77994
rect 4686 41758 4922 41994
rect 4686 5758 4922 5994
rect -3894 -2502 -3658 -2266
rect -3574 -2502 -3338 -2266
rect -3894 -2822 -3658 -2586
rect -3574 -2822 -3338 -2586
rect 4686 -2502 4922 -2266
rect 4686 -2822 4922 -2586
rect -4854 -3462 -4618 -3226
rect -4534 -3462 -4298 -3226
rect -4854 -3782 -4618 -3546
rect -4534 -3782 -4298 -3546
rect 8386 693458 8622 693694
rect 8386 657458 8622 657694
rect 8386 621458 8622 621694
rect 8386 585458 8622 585694
rect 8386 549458 8622 549694
rect 8386 513458 8622 513694
rect 8386 477458 8622 477694
rect 8386 441458 8622 441694
rect 8386 405458 8622 405694
rect 8386 369458 8622 369694
rect 8386 333458 8622 333694
rect 8386 297458 8622 297694
rect 8386 261458 8622 261694
rect 8386 225458 8622 225694
rect 8386 189458 8622 189694
rect 8386 153458 8622 153694
rect 8386 117458 8622 117694
rect 8386 81458 8622 81694
rect 8386 45458 8622 45694
rect 8386 9458 8622 9694
rect -5814 -4422 -5578 -4186
rect -5494 -4422 -5258 -4186
rect -5814 -4742 -5578 -4506
rect -5494 -4742 -5258 -4506
rect 8386 -4422 8622 -4186
rect 8386 -4742 8622 -4506
rect -6774 -5382 -6538 -5146
rect -6454 -5382 -6218 -5146
rect -6774 -5702 -6538 -5466
rect -6454 -5702 -6218 -5466
rect 30086 711322 30322 711558
rect 30086 711002 30322 711238
rect 26386 709402 26622 709638
rect 26386 709082 26622 709318
rect 22686 707482 22922 707718
rect 22686 707162 22922 707398
rect 12086 697158 12322 697394
rect 12086 661158 12322 661394
rect 12086 625158 12322 625394
rect 12086 589158 12322 589394
rect 12086 553158 12322 553394
rect 12086 517158 12322 517394
rect 12086 481158 12322 481394
rect 12086 445158 12322 445394
rect 12086 409158 12322 409394
rect 12086 373158 12322 373394
rect 12086 337158 12322 337394
rect 12086 301158 12322 301394
rect 12086 265158 12322 265394
rect 12086 229158 12322 229394
rect 12086 193158 12322 193394
rect 12086 157158 12322 157394
rect 12086 121158 12322 121394
rect 12086 85158 12322 85394
rect 12086 49158 12322 49394
rect 12086 13158 12322 13394
rect -7734 -6342 -7498 -6106
rect -7414 -6342 -7178 -6106
rect -7734 -6662 -7498 -6426
rect -7414 -6662 -7178 -6426
rect 18986 705562 19222 705798
rect 18986 705242 19222 705478
rect 18986 668058 19222 668294
rect 18986 632058 19222 632294
rect 18986 596058 19222 596294
rect 18986 560058 19222 560294
rect 18986 524058 19222 524294
rect 18986 488058 19222 488294
rect 18986 452058 19222 452294
rect 18986 416058 19222 416294
rect 18986 380058 19222 380294
rect 18986 344058 19222 344294
rect 18986 308058 19222 308294
rect 18986 272058 19222 272294
rect 18986 236058 19222 236294
rect 18986 200058 19222 200294
rect 18986 164058 19222 164294
rect 18986 128058 19222 128294
rect 18986 92058 19222 92294
rect 18986 56058 19222 56294
rect 18986 20058 19222 20294
rect 18986 -1542 19222 -1306
rect 18986 -1862 19222 -1626
rect 22686 671758 22922 671994
rect 22686 635758 22922 635994
rect 22686 599758 22922 599994
rect 22686 563758 22922 563994
rect 22686 527758 22922 527994
rect 22686 491758 22922 491994
rect 22686 455758 22922 455994
rect 22686 419758 22922 419994
rect 22686 383758 22922 383994
rect 22686 347758 22922 347994
rect 22686 311758 22922 311994
rect 22686 275758 22922 275994
rect 22686 239758 22922 239994
rect 22686 203758 22922 203994
rect 22686 167758 22922 167994
rect 22686 131758 22922 131994
rect 22686 95758 22922 95994
rect 22686 59758 22922 59994
rect 22686 23758 22922 23994
rect 22686 -3462 22922 -3226
rect 22686 -3782 22922 -3546
rect 26386 675458 26622 675694
rect 26386 639458 26622 639694
rect 26386 603458 26622 603694
rect 26386 567458 26622 567694
rect 26386 531458 26622 531694
rect 26386 495458 26622 495694
rect 26386 459458 26622 459694
rect 26386 423458 26622 423694
rect 26386 387458 26622 387694
rect 26386 351458 26622 351694
rect 26386 315458 26622 315694
rect 26386 279458 26622 279694
rect 26386 243458 26622 243694
rect 26386 207458 26622 207694
rect 26386 171458 26622 171694
rect 26386 135458 26622 135694
rect 26386 99458 26622 99694
rect 26386 63458 26622 63694
rect 26386 27458 26622 27694
rect 26386 -5382 26622 -5146
rect 26386 -5702 26622 -5466
rect 48086 710362 48322 710598
rect 48086 710042 48322 710278
rect 44386 708442 44622 708678
rect 44386 708122 44622 708358
rect 40686 706522 40922 706758
rect 40686 706202 40922 706438
rect 30086 679158 30322 679394
rect 30086 643158 30322 643394
rect 30086 607158 30322 607394
rect 30086 571158 30322 571394
rect 30086 535158 30322 535394
rect 30086 499158 30322 499394
rect 30086 463158 30322 463394
rect 30086 427158 30322 427394
rect 30086 391158 30322 391394
rect 30086 355158 30322 355394
rect 30086 319158 30322 319394
rect 30086 283158 30322 283394
rect 30086 247158 30322 247394
rect 30086 211158 30322 211394
rect 30086 175158 30322 175394
rect 30086 139158 30322 139394
rect 30086 103158 30322 103394
rect 30086 67158 30322 67394
rect 30086 31158 30322 31394
rect 12086 -6342 12322 -6106
rect 12086 -6662 12322 -6426
rect -8694 -7302 -8458 -7066
rect -8374 -7302 -8138 -7066
rect -8694 -7622 -8458 -7386
rect -8374 -7622 -8138 -7386
rect 36986 704602 37222 704838
rect 36986 704282 37222 704518
rect 36986 686058 37222 686294
rect 36986 650058 37222 650294
rect 36986 614058 37222 614294
rect 36986 578058 37222 578294
rect 36986 542058 37222 542294
rect 36986 506058 37222 506294
rect 36986 470058 37222 470294
rect 36986 434058 37222 434294
rect 40686 689758 40922 689994
rect 40686 653758 40922 653994
rect 40686 617758 40922 617994
rect 40686 581758 40922 581994
rect 40686 545758 40922 545994
rect 40686 509758 40922 509994
rect 40686 473758 40922 473994
rect 40686 437758 40922 437994
rect 44386 693458 44622 693694
rect 44386 657458 44622 657694
rect 44386 621458 44622 621694
rect 44386 585458 44622 585694
rect 44386 549458 44622 549694
rect 44386 513458 44622 513694
rect 44386 477458 44622 477694
rect 44386 441458 44622 441694
rect 66086 711322 66322 711558
rect 66086 711002 66322 711238
rect 62386 709402 62622 709638
rect 62386 709082 62622 709318
rect 58686 707482 58922 707718
rect 58686 707162 58922 707398
rect 48086 697158 48322 697394
rect 48086 661158 48322 661394
rect 48086 625158 48322 625394
rect 48086 589158 48322 589394
rect 48086 553158 48322 553394
rect 48086 517158 48322 517394
rect 48086 481158 48322 481394
rect 48086 445158 48322 445394
rect 54986 705562 55222 705798
rect 54986 705242 55222 705478
rect 54986 668058 55222 668294
rect 54986 632058 55222 632294
rect 54986 596058 55222 596294
rect 54986 560058 55222 560294
rect 54986 524058 55222 524294
rect 54986 488058 55222 488294
rect 54986 452058 55222 452294
rect 58686 671758 58922 671994
rect 58686 635758 58922 635994
rect 58686 599758 58922 599994
rect 58686 563758 58922 563994
rect 58686 527758 58922 527994
rect 58686 491758 58922 491994
rect 58686 455758 58922 455994
rect 62386 675458 62622 675694
rect 62386 639458 62622 639694
rect 62386 603458 62622 603694
rect 62386 567458 62622 567694
rect 62386 531458 62622 531694
rect 62386 495458 62622 495694
rect 62386 459458 62622 459694
rect 84086 710362 84322 710598
rect 84086 710042 84322 710278
rect 80386 708442 80622 708678
rect 80386 708122 80622 708358
rect 76686 706522 76922 706758
rect 76686 706202 76922 706438
rect 66086 679158 66322 679394
rect 66086 643158 66322 643394
rect 66086 607158 66322 607394
rect 66086 571158 66322 571394
rect 66086 535158 66322 535394
rect 66086 499158 66322 499394
rect 66086 463158 66322 463394
rect 66086 427158 66322 427394
rect 72986 704602 73222 704838
rect 72986 704282 73222 704518
rect 72986 686058 73222 686294
rect 72986 650058 73222 650294
rect 72986 614058 73222 614294
rect 72986 578058 73222 578294
rect 72986 542058 73222 542294
rect 72986 506058 73222 506294
rect 72986 470058 73222 470294
rect 72986 434058 73222 434294
rect 76686 689758 76922 689994
rect 76686 653758 76922 653994
rect 76686 617758 76922 617994
rect 76686 581758 76922 581994
rect 76686 545758 76922 545994
rect 76686 509758 76922 509994
rect 76686 473758 76922 473994
rect 76686 437758 76922 437994
rect 80386 693458 80622 693694
rect 80386 657458 80622 657694
rect 80386 621458 80622 621694
rect 80386 585458 80622 585694
rect 80386 549458 80622 549694
rect 80386 513458 80622 513694
rect 80386 477458 80622 477694
rect 80386 441458 80622 441694
rect 102086 711322 102322 711558
rect 102086 711002 102322 711238
rect 98386 709402 98622 709638
rect 98386 709082 98622 709318
rect 94686 707482 94922 707718
rect 94686 707162 94922 707398
rect 84086 697158 84322 697394
rect 84086 661158 84322 661394
rect 84086 625158 84322 625394
rect 84086 589158 84322 589394
rect 84086 553158 84322 553394
rect 84086 517158 84322 517394
rect 84086 481158 84322 481394
rect 84086 445158 84322 445394
rect 90986 705562 91222 705798
rect 90986 705242 91222 705478
rect 90986 668058 91222 668294
rect 90986 632058 91222 632294
rect 90986 596058 91222 596294
rect 90986 560058 91222 560294
rect 90986 524058 91222 524294
rect 90986 488058 91222 488294
rect 90986 452058 91222 452294
rect 94686 671758 94922 671994
rect 94686 635758 94922 635994
rect 94686 599758 94922 599994
rect 94686 563758 94922 563994
rect 94686 527758 94922 527994
rect 94686 491758 94922 491994
rect 94686 455758 94922 455994
rect 98386 675458 98622 675694
rect 98386 639458 98622 639694
rect 98386 603458 98622 603694
rect 98386 567458 98622 567694
rect 98386 531458 98622 531694
rect 98386 495458 98622 495694
rect 98386 459458 98622 459694
rect 120086 710362 120322 710598
rect 120086 710042 120322 710278
rect 116386 708442 116622 708678
rect 116386 708122 116622 708358
rect 112686 706522 112922 706758
rect 112686 706202 112922 706438
rect 102086 679158 102322 679394
rect 102086 643158 102322 643394
rect 102086 607158 102322 607394
rect 102086 571158 102322 571394
rect 102086 535158 102322 535394
rect 102086 499158 102322 499394
rect 102086 463158 102322 463394
rect 102086 427158 102322 427394
rect 108986 704602 109222 704838
rect 108986 704282 109222 704518
rect 108986 686058 109222 686294
rect 108986 650058 109222 650294
rect 108986 614058 109222 614294
rect 108986 578058 109222 578294
rect 108986 542058 109222 542294
rect 108986 506058 109222 506294
rect 108986 470058 109222 470294
rect 108986 434058 109222 434294
rect 112686 689758 112922 689994
rect 112686 653758 112922 653994
rect 112686 617758 112922 617994
rect 112686 581758 112922 581994
rect 112686 545758 112922 545994
rect 112686 509758 112922 509994
rect 112686 473758 112922 473994
rect 112686 437758 112922 437994
rect 116386 693458 116622 693694
rect 116386 657458 116622 657694
rect 116386 621458 116622 621694
rect 116386 585458 116622 585694
rect 116386 549458 116622 549694
rect 116386 513458 116622 513694
rect 116386 477458 116622 477694
rect 116386 441458 116622 441694
rect 138086 711322 138322 711558
rect 138086 711002 138322 711238
rect 134386 709402 134622 709638
rect 134386 709082 134622 709318
rect 130686 707482 130922 707718
rect 130686 707162 130922 707398
rect 120086 697158 120322 697394
rect 120086 661158 120322 661394
rect 120086 625158 120322 625394
rect 120086 589158 120322 589394
rect 120086 553158 120322 553394
rect 120086 517158 120322 517394
rect 120086 481158 120322 481394
rect 120086 445158 120322 445394
rect 126986 705562 127222 705798
rect 126986 705242 127222 705478
rect 126986 668058 127222 668294
rect 126986 632058 127222 632294
rect 126986 596058 127222 596294
rect 126986 560058 127222 560294
rect 126986 524058 127222 524294
rect 126986 488058 127222 488294
rect 126986 452058 127222 452294
rect 130686 671758 130922 671994
rect 130686 635758 130922 635994
rect 130686 599758 130922 599994
rect 130686 563758 130922 563994
rect 130686 527758 130922 527994
rect 130686 491758 130922 491994
rect 130686 455758 130922 455994
rect 134386 675458 134622 675694
rect 134386 639458 134622 639694
rect 134386 603458 134622 603694
rect 134386 567458 134622 567694
rect 134386 531458 134622 531694
rect 134386 495458 134622 495694
rect 134386 459458 134622 459694
rect 156086 710362 156322 710598
rect 156086 710042 156322 710278
rect 152386 708442 152622 708678
rect 152386 708122 152622 708358
rect 148686 706522 148922 706758
rect 148686 706202 148922 706438
rect 138086 679158 138322 679394
rect 138086 643158 138322 643394
rect 138086 607158 138322 607394
rect 138086 571158 138322 571394
rect 138086 535158 138322 535394
rect 138086 499158 138322 499394
rect 138086 463158 138322 463394
rect 138086 427158 138322 427394
rect 144986 704602 145222 704838
rect 144986 704282 145222 704518
rect 144986 686058 145222 686294
rect 144986 650058 145222 650294
rect 144986 614058 145222 614294
rect 144986 578058 145222 578294
rect 144986 542058 145222 542294
rect 144986 506058 145222 506294
rect 144986 470058 145222 470294
rect 144986 434058 145222 434294
rect 148686 689758 148922 689994
rect 148686 653758 148922 653994
rect 148686 617758 148922 617994
rect 148686 581758 148922 581994
rect 148686 545758 148922 545994
rect 148686 509758 148922 509994
rect 148686 473758 148922 473994
rect 148686 437758 148922 437994
rect 152386 693458 152622 693694
rect 152386 657458 152622 657694
rect 152386 621458 152622 621694
rect 152386 585458 152622 585694
rect 152386 549458 152622 549694
rect 152386 513458 152622 513694
rect 152386 477458 152622 477694
rect 152386 441458 152622 441694
rect 174086 711322 174322 711558
rect 174086 711002 174322 711238
rect 170386 709402 170622 709638
rect 170386 709082 170622 709318
rect 166686 707482 166922 707718
rect 166686 707162 166922 707398
rect 156086 697158 156322 697394
rect 156086 661158 156322 661394
rect 156086 625158 156322 625394
rect 156086 589158 156322 589394
rect 156086 553158 156322 553394
rect 156086 517158 156322 517394
rect 156086 481158 156322 481394
rect 156086 445158 156322 445394
rect 162986 705562 163222 705798
rect 162986 705242 163222 705478
rect 162986 668058 163222 668294
rect 162986 632058 163222 632294
rect 162986 596058 163222 596294
rect 162986 560058 163222 560294
rect 162986 524058 163222 524294
rect 162986 488058 163222 488294
rect 162986 452058 163222 452294
rect 166686 671758 166922 671994
rect 166686 635758 166922 635994
rect 166686 599758 166922 599994
rect 166686 563758 166922 563994
rect 166686 527758 166922 527994
rect 166686 491758 166922 491994
rect 166686 455758 166922 455994
rect 170386 675458 170622 675694
rect 170386 639458 170622 639694
rect 170386 603458 170622 603694
rect 170386 567458 170622 567694
rect 170386 531458 170622 531694
rect 170386 495458 170622 495694
rect 170386 459458 170622 459694
rect 192086 710362 192322 710598
rect 192086 710042 192322 710278
rect 188386 708442 188622 708678
rect 188386 708122 188622 708358
rect 184686 706522 184922 706758
rect 184686 706202 184922 706438
rect 174086 679158 174322 679394
rect 174086 643158 174322 643394
rect 174086 607158 174322 607394
rect 174086 571158 174322 571394
rect 174086 535158 174322 535394
rect 174086 499158 174322 499394
rect 174086 463158 174322 463394
rect 174086 427158 174322 427394
rect 180986 704602 181222 704838
rect 180986 704282 181222 704518
rect 180986 686058 181222 686294
rect 180986 650058 181222 650294
rect 180986 614058 181222 614294
rect 180986 578058 181222 578294
rect 180986 542058 181222 542294
rect 180986 506058 181222 506294
rect 180986 470058 181222 470294
rect 180986 434058 181222 434294
rect 40328 416058 40564 416294
rect 176056 416058 176292 416294
rect 36986 398058 37222 398294
rect 41008 398058 41244 398294
rect 175376 398058 175612 398294
rect 180986 398058 181222 398294
rect 40328 380058 40564 380294
rect 176056 380058 176292 380294
rect 36986 362058 37222 362294
rect 41008 362058 41244 362294
rect 175376 362058 175612 362294
rect 180986 362058 181222 362294
rect 40328 344058 40564 344294
rect 176056 344058 176292 344294
rect 36986 326058 37222 326294
rect 36986 290058 37222 290294
rect 36986 254058 37222 254294
rect 40686 329758 40922 329994
rect 40686 293758 40922 293994
rect 40686 257758 40922 257994
rect 44386 333458 44622 333694
rect 44386 297458 44622 297694
rect 44386 261458 44622 261694
rect 48086 337158 48322 337394
rect 48086 301158 48322 301394
rect 48086 265158 48322 265394
rect 36986 218058 37222 218294
rect 44250 218058 44486 218294
rect 36986 182058 37222 182294
rect 44250 182058 44486 182294
rect 36986 146058 37222 146294
rect 44250 146058 44486 146294
rect 36986 110058 37222 110294
rect 44250 110058 44486 110294
rect 36986 74058 37222 74294
rect 44250 74058 44486 74294
rect 36986 38058 37222 38294
rect 36986 2058 37222 2294
rect 36986 -582 37222 -346
rect 36986 -902 37222 -666
rect 40686 5758 40922 5994
rect 40686 -2502 40922 -2266
rect 40686 -2822 40922 -2586
rect 44386 9458 44622 9694
rect 44386 -4422 44622 -4186
rect 44386 -4742 44622 -4506
rect 54986 308058 55222 308294
rect 54986 272058 55222 272294
rect 48086 13158 48322 13394
rect 30086 -7302 30322 -7066
rect 30086 -7622 30322 -7386
rect 58686 311758 58922 311994
rect 58686 275758 58922 275994
rect 62386 315458 62622 315694
rect 62386 279458 62622 279694
rect 62386 243458 62622 243694
rect 66086 319158 66322 319394
rect 66086 283158 66322 283394
rect 66086 247158 66322 247394
rect 72986 326058 73222 326294
rect 72986 290058 73222 290294
rect 72986 254058 73222 254294
rect 76686 329758 76922 329994
rect 76686 293758 76922 293994
rect 76686 257758 76922 257994
rect 80386 333458 80622 333694
rect 80386 297458 80622 297694
rect 80386 261458 80622 261694
rect 84086 337158 84322 337394
rect 84086 301158 84322 301394
rect 84086 265158 84322 265394
rect 90986 308058 91222 308294
rect 90986 272058 91222 272294
rect 94686 311758 94922 311994
rect 94686 275758 94922 275994
rect 98386 315458 98622 315694
rect 98386 279458 98622 279694
rect 98386 243458 98622 243694
rect 102086 319158 102322 319394
rect 102086 283158 102322 283394
rect 102086 247158 102322 247394
rect 108986 326058 109222 326294
rect 108986 290058 109222 290294
rect 108986 254058 109222 254294
rect 112686 329758 112922 329994
rect 112686 293758 112922 293994
rect 112686 257758 112922 257994
rect 116386 333458 116622 333694
rect 116386 297458 116622 297694
rect 116386 261458 116622 261694
rect 120086 337158 120322 337394
rect 120086 301158 120322 301394
rect 120086 265158 120322 265394
rect 126986 308058 127222 308294
rect 126986 272058 127222 272294
rect 130686 311758 130922 311994
rect 130686 275758 130922 275994
rect 134386 315458 134622 315694
rect 134386 279458 134622 279694
rect 134386 243458 134622 243694
rect 138086 319158 138322 319394
rect 138086 283158 138322 283394
rect 138086 247158 138322 247394
rect 144986 326058 145222 326294
rect 144986 290058 145222 290294
rect 144986 254058 145222 254294
rect 148686 329758 148922 329994
rect 148686 293758 148922 293994
rect 148686 257758 148922 257994
rect 152386 333458 152622 333694
rect 152386 297458 152622 297694
rect 152386 261458 152622 261694
rect 156086 337158 156322 337394
rect 156086 301158 156322 301394
rect 156086 265158 156322 265394
rect 162986 308058 163222 308294
rect 162986 272058 163222 272294
rect 166686 311758 166922 311994
rect 166686 275758 166922 275994
rect 170386 315458 170622 315694
rect 170386 279458 170622 279694
rect 170386 243458 170622 243694
rect 174086 319158 174322 319394
rect 174086 283158 174322 283394
rect 174086 247158 174322 247394
rect 180986 326058 181222 326294
rect 180986 290058 181222 290294
rect 180986 254058 181222 254294
rect 184686 689758 184922 689994
rect 184686 653758 184922 653994
rect 184686 617758 184922 617994
rect 184686 581758 184922 581994
rect 184686 545758 184922 545994
rect 184686 509758 184922 509994
rect 184686 473758 184922 473994
rect 184686 437758 184922 437994
rect 184686 401758 184922 401994
rect 184686 365758 184922 365994
rect 184686 329758 184922 329994
rect 184686 293758 184922 293994
rect 184686 257758 184922 257994
rect 188386 693458 188622 693694
rect 188386 657458 188622 657694
rect 188386 621458 188622 621694
rect 188386 585458 188622 585694
rect 188386 549458 188622 549694
rect 188386 513458 188622 513694
rect 188386 477458 188622 477694
rect 188386 441458 188622 441694
rect 188386 405458 188622 405694
rect 188386 369458 188622 369694
rect 188386 333458 188622 333694
rect 188386 297458 188622 297694
rect 188386 261458 188622 261694
rect 210086 711322 210322 711558
rect 210086 711002 210322 711238
rect 206386 709402 206622 709638
rect 206386 709082 206622 709318
rect 202686 707482 202922 707718
rect 202686 707162 202922 707398
rect 192086 697158 192322 697394
rect 192086 661158 192322 661394
rect 192086 625158 192322 625394
rect 192086 589158 192322 589394
rect 192086 553158 192322 553394
rect 192086 517158 192322 517394
rect 192086 481158 192322 481394
rect 192086 445158 192322 445394
rect 192086 409158 192322 409394
rect 192086 373158 192322 373394
rect 192086 337158 192322 337394
rect 192086 301158 192322 301394
rect 192086 265158 192322 265394
rect 198986 705562 199222 705798
rect 198986 705242 199222 705478
rect 198986 668058 199222 668294
rect 198986 632058 199222 632294
rect 198986 596058 199222 596294
rect 198986 560058 199222 560294
rect 198986 524058 199222 524294
rect 198986 488058 199222 488294
rect 198986 452058 199222 452294
rect 198986 416058 199222 416294
rect 198986 380058 199222 380294
rect 198986 344058 199222 344294
rect 198986 308058 199222 308294
rect 198986 272058 199222 272294
rect 202686 671758 202922 671994
rect 202686 635758 202922 635994
rect 202686 599758 202922 599994
rect 202686 563758 202922 563994
rect 202686 527758 202922 527994
rect 202686 491758 202922 491994
rect 202686 455758 202922 455994
rect 202686 419758 202922 419994
rect 202686 383758 202922 383994
rect 202686 347758 202922 347994
rect 202686 311758 202922 311994
rect 202686 275758 202922 275994
rect 206386 675458 206622 675694
rect 206386 639458 206622 639694
rect 206386 603458 206622 603694
rect 206386 567458 206622 567694
rect 206386 531458 206622 531694
rect 206386 495458 206622 495694
rect 206386 459458 206622 459694
rect 206386 423458 206622 423694
rect 206386 387458 206622 387694
rect 206386 351458 206622 351694
rect 206386 315458 206622 315694
rect 206386 279458 206622 279694
rect 206386 243458 206622 243694
rect 228086 710362 228322 710598
rect 228086 710042 228322 710278
rect 224386 708442 224622 708678
rect 224386 708122 224622 708358
rect 220686 706522 220922 706758
rect 220686 706202 220922 706438
rect 210086 679158 210322 679394
rect 210086 643158 210322 643394
rect 210086 607158 210322 607394
rect 210086 571158 210322 571394
rect 210086 535158 210322 535394
rect 210086 499158 210322 499394
rect 210086 463158 210322 463394
rect 210086 427158 210322 427394
rect 210086 391158 210322 391394
rect 210086 355158 210322 355394
rect 210086 319158 210322 319394
rect 210086 283158 210322 283394
rect 210086 247158 210322 247394
rect 216986 704602 217222 704838
rect 216986 704282 217222 704518
rect 216986 686058 217222 686294
rect 216986 650058 217222 650294
rect 216986 614058 217222 614294
rect 216986 578058 217222 578294
rect 216986 542058 217222 542294
rect 216986 506058 217222 506294
rect 216986 470058 217222 470294
rect 216986 434058 217222 434294
rect 216986 398058 217222 398294
rect 216986 362058 217222 362294
rect 216986 326058 217222 326294
rect 216986 290058 217222 290294
rect 216986 254058 217222 254294
rect 220686 689758 220922 689994
rect 220686 653758 220922 653994
rect 220686 617758 220922 617994
rect 220686 581758 220922 581994
rect 220686 545758 220922 545994
rect 220686 509758 220922 509994
rect 220686 473758 220922 473994
rect 220686 437758 220922 437994
rect 220686 401758 220922 401994
rect 220686 365758 220922 365994
rect 220686 329758 220922 329994
rect 220686 293758 220922 293994
rect 220686 257758 220922 257994
rect 224386 693458 224622 693694
rect 224386 657458 224622 657694
rect 224386 621458 224622 621694
rect 224386 585458 224622 585694
rect 224386 549458 224622 549694
rect 224386 513458 224622 513694
rect 224386 477458 224622 477694
rect 224386 441458 224622 441694
rect 224386 405458 224622 405694
rect 224386 369458 224622 369694
rect 224386 333458 224622 333694
rect 224386 297458 224622 297694
rect 224386 261458 224622 261694
rect 246086 711322 246322 711558
rect 246086 711002 246322 711238
rect 242386 709402 242622 709638
rect 242386 709082 242622 709318
rect 238686 707482 238922 707718
rect 238686 707162 238922 707398
rect 228086 697158 228322 697394
rect 228086 661158 228322 661394
rect 228086 625158 228322 625394
rect 228086 589158 228322 589394
rect 228086 553158 228322 553394
rect 228086 517158 228322 517394
rect 228086 481158 228322 481394
rect 228086 445158 228322 445394
rect 228086 409158 228322 409394
rect 228086 373158 228322 373394
rect 234986 705562 235222 705798
rect 234986 705242 235222 705478
rect 234986 668058 235222 668294
rect 234986 632058 235222 632294
rect 234986 596058 235222 596294
rect 234986 560058 235222 560294
rect 234986 524058 235222 524294
rect 234986 488058 235222 488294
rect 234986 452058 235222 452294
rect 234986 416058 235222 416294
rect 234986 380058 235222 380294
rect 234986 344058 235222 344294
rect 228086 337158 228322 337394
rect 228086 301158 228322 301394
rect 228086 265158 228322 265394
rect 59610 236058 59846 236294
rect 90330 236058 90566 236294
rect 121050 236058 121286 236294
rect 151770 236058 152006 236294
rect 182490 236058 182726 236294
rect 213210 236058 213446 236294
rect 74970 218058 75206 218294
rect 105690 218058 105926 218294
rect 136410 218058 136646 218294
rect 167130 218058 167366 218294
rect 197850 218058 198086 218294
rect 228570 218058 228806 218294
rect 59610 200058 59846 200294
rect 90330 200058 90566 200294
rect 121050 200058 121286 200294
rect 151770 200058 152006 200294
rect 182490 200058 182726 200294
rect 213210 200058 213446 200294
rect 74970 182058 75206 182294
rect 105690 182058 105926 182294
rect 136410 182058 136646 182294
rect 167130 182058 167366 182294
rect 197850 182058 198086 182294
rect 228570 182058 228806 182294
rect 59610 164058 59846 164294
rect 90330 164058 90566 164294
rect 121050 164058 121286 164294
rect 151770 164058 152006 164294
rect 182490 164058 182726 164294
rect 213210 164058 213446 164294
rect 74970 146058 75206 146294
rect 105690 146058 105926 146294
rect 136410 146058 136646 146294
rect 167130 146058 167366 146294
rect 197850 146058 198086 146294
rect 228570 146058 228806 146294
rect 59610 128058 59846 128294
rect 90330 128058 90566 128294
rect 121050 128058 121286 128294
rect 151770 128058 152006 128294
rect 182490 128058 182726 128294
rect 213210 128058 213446 128294
rect 74970 110058 75206 110294
rect 105690 110058 105926 110294
rect 136410 110058 136646 110294
rect 167130 110058 167366 110294
rect 197850 110058 198086 110294
rect 228570 110058 228806 110294
rect 59610 92058 59846 92294
rect 90330 92058 90566 92294
rect 121050 92058 121286 92294
rect 151770 92058 152006 92294
rect 182490 92058 182726 92294
rect 213210 92058 213446 92294
rect 74970 74058 75206 74294
rect 105690 74058 105926 74294
rect 136410 74058 136646 74294
rect 167130 74058 167366 74294
rect 197850 74058 198086 74294
rect 228570 74058 228806 74294
rect 59610 56058 59846 56294
rect 90330 56058 90566 56294
rect 121050 56058 121286 56294
rect 151770 56058 152006 56294
rect 182490 56058 182726 56294
rect 213210 56058 213446 56294
rect 234986 308058 235222 308294
rect 234986 272058 235222 272294
rect 238686 671758 238922 671994
rect 238686 635758 238922 635994
rect 238686 599758 238922 599994
rect 238686 563758 238922 563994
rect 238686 527758 238922 527994
rect 238686 491758 238922 491994
rect 238686 455758 238922 455994
rect 238686 419758 238922 419994
rect 238686 383758 238922 383994
rect 238686 347758 238922 347994
rect 238686 311758 238922 311994
rect 238686 275758 238922 275994
rect 242386 675458 242622 675694
rect 242386 639458 242622 639694
rect 242386 603458 242622 603694
rect 242386 567458 242622 567694
rect 242386 531458 242622 531694
rect 242386 495458 242622 495694
rect 242386 459458 242622 459694
rect 242386 423458 242622 423694
rect 242386 387458 242622 387694
rect 242386 351458 242622 351694
rect 242386 315458 242622 315694
rect 242386 279458 242622 279694
rect 242386 243458 242622 243694
rect 242386 207458 242622 207694
rect 242386 171458 242622 171694
rect 242386 135458 242622 135694
rect 242386 99458 242622 99694
rect 242386 63458 242622 63694
rect 54986 20058 55222 20294
rect 54986 -1542 55222 -1306
rect 54986 -1862 55222 -1626
rect 58686 23758 58922 23994
rect 58686 -3462 58922 -3226
rect 58686 -3782 58922 -3546
rect 62386 27458 62622 27694
rect 62386 -5382 62622 -5146
rect 62386 -5702 62622 -5466
rect 66086 31158 66322 31394
rect 48086 -6342 48322 -6106
rect 48086 -6662 48322 -6426
rect 72986 2058 73222 2294
rect 72986 -582 73222 -346
rect 72986 -902 73222 -666
rect 76686 5758 76922 5994
rect 76686 -2502 76922 -2266
rect 76686 -2822 76922 -2586
rect 80386 9458 80622 9694
rect 80386 -4422 80622 -4186
rect 80386 -4742 80622 -4506
rect 84086 13158 84322 13394
rect 66086 -7302 66322 -7066
rect 66086 -7622 66322 -7386
rect 90986 20058 91222 20294
rect 90986 -1542 91222 -1306
rect 90986 -1862 91222 -1626
rect 94686 23758 94922 23994
rect 94686 -3462 94922 -3226
rect 94686 -3782 94922 -3546
rect 98386 27458 98622 27694
rect 98386 -5382 98622 -5146
rect 98386 -5702 98622 -5466
rect 102086 31158 102322 31394
rect 84086 -6342 84322 -6106
rect 84086 -6662 84322 -6426
rect 108986 2058 109222 2294
rect 108986 -582 109222 -346
rect 108986 -902 109222 -666
rect 112686 5758 112922 5994
rect 112686 -2502 112922 -2266
rect 112686 -2822 112922 -2586
rect 116386 9458 116622 9694
rect 116386 -4422 116622 -4186
rect 116386 -4742 116622 -4506
rect 120086 13158 120322 13394
rect 102086 -7302 102322 -7066
rect 102086 -7622 102322 -7386
rect 126986 20058 127222 20294
rect 126986 -1542 127222 -1306
rect 126986 -1862 127222 -1626
rect 130686 23758 130922 23994
rect 130686 -3462 130922 -3226
rect 130686 -3782 130922 -3546
rect 134386 27458 134622 27694
rect 134386 -5382 134622 -5146
rect 134386 -5702 134622 -5466
rect 138086 31158 138322 31394
rect 120086 -6342 120322 -6106
rect 120086 -6662 120322 -6426
rect 144986 2058 145222 2294
rect 144986 -582 145222 -346
rect 144986 -902 145222 -666
rect 148686 5758 148922 5994
rect 148686 -2502 148922 -2266
rect 148686 -2822 148922 -2586
rect 152386 9458 152622 9694
rect 152386 -4422 152622 -4186
rect 152386 -4742 152622 -4506
rect 156086 13158 156322 13394
rect 138086 -7302 138322 -7066
rect 138086 -7622 138322 -7386
rect 162986 20058 163222 20294
rect 162986 -1542 163222 -1306
rect 162986 -1862 163222 -1626
rect 166686 23758 166922 23994
rect 166686 -3462 166922 -3226
rect 166686 -3782 166922 -3546
rect 170386 27458 170622 27694
rect 170386 -5382 170622 -5146
rect 170386 -5702 170622 -5466
rect 174086 31158 174322 31394
rect 156086 -6342 156322 -6106
rect 156086 -6662 156322 -6426
rect 180986 2058 181222 2294
rect 180986 -582 181222 -346
rect 180986 -902 181222 -666
rect 184686 5758 184922 5994
rect 184686 -2502 184922 -2266
rect 184686 -2822 184922 -2586
rect 188386 9458 188622 9694
rect 188386 -4422 188622 -4186
rect 188386 -4742 188622 -4506
rect 192086 13158 192322 13394
rect 174086 -7302 174322 -7066
rect 174086 -7622 174322 -7386
rect 198986 20058 199222 20294
rect 198986 -1542 199222 -1306
rect 198986 -1862 199222 -1626
rect 202686 23758 202922 23994
rect 202686 -3462 202922 -3226
rect 202686 -3782 202922 -3546
rect 206386 27458 206622 27694
rect 206386 -5382 206622 -5146
rect 206386 -5702 206622 -5466
rect 210086 31158 210322 31394
rect 192086 -6342 192322 -6106
rect 192086 -6662 192322 -6426
rect 216986 2058 217222 2294
rect 216986 -582 217222 -346
rect 216986 -902 217222 -666
rect 220686 5758 220922 5994
rect 220686 -2502 220922 -2266
rect 220686 -2822 220922 -2586
rect 224386 9458 224622 9694
rect 224386 -4422 224622 -4186
rect 224386 -4742 224622 -4506
rect 228086 13158 228322 13394
rect 210086 -7302 210322 -7066
rect 210086 -7622 210322 -7386
rect 234986 20058 235222 20294
rect 234986 -1542 235222 -1306
rect 234986 -1862 235222 -1626
rect 238686 23758 238922 23994
rect 238686 -3462 238922 -3226
rect 238686 -3782 238922 -3546
rect 242386 27458 242622 27694
rect 242386 -5382 242622 -5146
rect 242386 -5702 242622 -5466
rect 264086 710362 264322 710598
rect 264086 710042 264322 710278
rect 260386 708442 260622 708678
rect 260386 708122 260622 708358
rect 256686 706522 256922 706758
rect 256686 706202 256922 706438
rect 246086 679158 246322 679394
rect 246086 643158 246322 643394
rect 246086 607158 246322 607394
rect 246086 571158 246322 571394
rect 246086 535158 246322 535394
rect 246086 499158 246322 499394
rect 246086 463158 246322 463394
rect 246086 427158 246322 427394
rect 246086 391158 246322 391394
rect 246086 355158 246322 355394
rect 246086 319158 246322 319394
rect 246086 283158 246322 283394
rect 246086 247158 246322 247394
rect 246086 211158 246322 211394
rect 246086 175158 246322 175394
rect 246086 139158 246322 139394
rect 246086 103158 246322 103394
rect 246086 67158 246322 67394
rect 246086 31158 246322 31394
rect 228086 -6342 228322 -6106
rect 228086 -6662 228322 -6426
rect 252986 704602 253222 704838
rect 252986 704282 253222 704518
rect 252986 686058 253222 686294
rect 252986 650058 253222 650294
rect 252986 614058 253222 614294
rect 252986 578058 253222 578294
rect 252986 542058 253222 542294
rect 252986 506058 253222 506294
rect 252986 470058 253222 470294
rect 252986 434058 253222 434294
rect 252986 398058 253222 398294
rect 252986 362058 253222 362294
rect 252986 326058 253222 326294
rect 252986 290058 253222 290294
rect 252986 254058 253222 254294
rect 252986 218058 253222 218294
rect 252986 182058 253222 182294
rect 252986 146058 253222 146294
rect 252986 110058 253222 110294
rect 252986 74058 253222 74294
rect 252986 38058 253222 38294
rect 252986 2058 253222 2294
rect 252986 -582 253222 -346
rect 252986 -902 253222 -666
rect 256686 689758 256922 689994
rect 256686 653758 256922 653994
rect 256686 617758 256922 617994
rect 256686 581758 256922 581994
rect 256686 545758 256922 545994
rect 256686 509758 256922 509994
rect 256686 473758 256922 473994
rect 256686 437758 256922 437994
rect 256686 401758 256922 401994
rect 256686 365758 256922 365994
rect 256686 329758 256922 329994
rect 256686 293758 256922 293994
rect 256686 257758 256922 257994
rect 256686 221758 256922 221994
rect 256686 185758 256922 185994
rect 256686 149758 256922 149994
rect 256686 113758 256922 113994
rect 256686 77758 256922 77994
rect 256686 41758 256922 41994
rect 256686 5758 256922 5994
rect 256686 -2502 256922 -2266
rect 256686 -2822 256922 -2586
rect 260386 693458 260622 693694
rect 260386 657458 260622 657694
rect 260386 621458 260622 621694
rect 260386 585458 260622 585694
rect 260386 549458 260622 549694
rect 260386 513458 260622 513694
rect 260386 477458 260622 477694
rect 260386 441458 260622 441694
rect 260386 405458 260622 405694
rect 260386 369458 260622 369694
rect 260386 333458 260622 333694
rect 260386 297458 260622 297694
rect 260386 261458 260622 261694
rect 260386 225458 260622 225694
rect 260386 189458 260622 189694
rect 260386 153458 260622 153694
rect 260386 117458 260622 117694
rect 260386 81458 260622 81694
rect 260386 45458 260622 45694
rect 260386 9458 260622 9694
rect 260386 -4422 260622 -4186
rect 260386 -4742 260622 -4506
rect 282086 711322 282322 711558
rect 282086 711002 282322 711238
rect 278386 709402 278622 709638
rect 278386 709082 278622 709318
rect 274686 707482 274922 707718
rect 274686 707162 274922 707398
rect 264086 697158 264322 697394
rect 264086 661158 264322 661394
rect 264086 625158 264322 625394
rect 264086 589158 264322 589394
rect 264086 553158 264322 553394
rect 264086 517158 264322 517394
rect 264086 481158 264322 481394
rect 264086 445158 264322 445394
rect 264086 409158 264322 409394
rect 264086 373158 264322 373394
rect 264086 337158 264322 337394
rect 264086 301158 264322 301394
rect 264086 265158 264322 265394
rect 264086 229158 264322 229394
rect 264086 193158 264322 193394
rect 264086 157158 264322 157394
rect 264086 121158 264322 121394
rect 264086 85158 264322 85394
rect 264086 49158 264322 49394
rect 264086 13158 264322 13394
rect 246086 -7302 246322 -7066
rect 246086 -7622 246322 -7386
rect 270986 705562 271222 705798
rect 270986 705242 271222 705478
rect 270986 668058 271222 668294
rect 270986 632058 271222 632294
rect 270986 596058 271222 596294
rect 270986 560058 271222 560294
rect 270986 524058 271222 524294
rect 270986 488058 271222 488294
rect 270986 452058 271222 452294
rect 270986 416058 271222 416294
rect 270986 380058 271222 380294
rect 270986 344058 271222 344294
rect 270986 308058 271222 308294
rect 270986 272058 271222 272294
rect 270986 236058 271222 236294
rect 270986 200058 271222 200294
rect 270986 164058 271222 164294
rect 270986 128058 271222 128294
rect 270986 92058 271222 92294
rect 270986 56058 271222 56294
rect 270986 20058 271222 20294
rect 270986 -1542 271222 -1306
rect 270986 -1862 271222 -1626
rect 274686 671758 274922 671994
rect 274686 635758 274922 635994
rect 274686 599758 274922 599994
rect 274686 563758 274922 563994
rect 274686 527758 274922 527994
rect 274686 491758 274922 491994
rect 274686 455758 274922 455994
rect 274686 419758 274922 419994
rect 274686 383758 274922 383994
rect 274686 347758 274922 347994
rect 274686 311758 274922 311994
rect 274686 275758 274922 275994
rect 274686 239758 274922 239994
rect 274686 203758 274922 203994
rect 274686 167758 274922 167994
rect 274686 131758 274922 131994
rect 274686 95758 274922 95994
rect 274686 59758 274922 59994
rect 274686 23758 274922 23994
rect 274686 -3462 274922 -3226
rect 274686 -3782 274922 -3546
rect 278386 675458 278622 675694
rect 278386 639458 278622 639694
rect 278386 603458 278622 603694
rect 278386 567458 278622 567694
rect 278386 531458 278622 531694
rect 278386 495458 278622 495694
rect 278386 459458 278622 459694
rect 278386 423458 278622 423694
rect 278386 387458 278622 387694
rect 278386 351458 278622 351694
rect 278386 315458 278622 315694
rect 278386 279458 278622 279694
rect 278386 243458 278622 243694
rect 278386 207458 278622 207694
rect 278386 171458 278622 171694
rect 278386 135458 278622 135694
rect 278386 99458 278622 99694
rect 278386 63458 278622 63694
rect 278386 27458 278622 27694
rect 278386 -5382 278622 -5146
rect 278386 -5702 278622 -5466
rect 300086 710362 300322 710598
rect 300086 710042 300322 710278
rect 296386 708442 296622 708678
rect 296386 708122 296622 708358
rect 292686 706522 292922 706758
rect 292686 706202 292922 706438
rect 282086 679158 282322 679394
rect 282086 643158 282322 643394
rect 282086 607158 282322 607394
rect 282086 571158 282322 571394
rect 282086 535158 282322 535394
rect 282086 499158 282322 499394
rect 282086 463158 282322 463394
rect 282086 427158 282322 427394
rect 282086 391158 282322 391394
rect 282086 355158 282322 355394
rect 282086 319158 282322 319394
rect 282086 283158 282322 283394
rect 282086 247158 282322 247394
rect 282086 211158 282322 211394
rect 282086 175158 282322 175394
rect 282086 139158 282322 139394
rect 282086 103158 282322 103394
rect 282086 67158 282322 67394
rect 282086 31158 282322 31394
rect 264086 -6342 264322 -6106
rect 264086 -6662 264322 -6426
rect 288986 704602 289222 704838
rect 288986 704282 289222 704518
rect 288986 686058 289222 686294
rect 288986 650058 289222 650294
rect 288986 614058 289222 614294
rect 288986 578058 289222 578294
rect 288986 542058 289222 542294
rect 288986 506058 289222 506294
rect 288986 470058 289222 470294
rect 288986 434058 289222 434294
rect 288986 398058 289222 398294
rect 288986 362058 289222 362294
rect 288986 326058 289222 326294
rect 288986 290058 289222 290294
rect 288986 254058 289222 254294
rect 288986 218058 289222 218294
rect 288986 182058 289222 182294
rect 288986 146058 289222 146294
rect 288986 110058 289222 110294
rect 288986 74058 289222 74294
rect 288986 38058 289222 38294
rect 288986 2058 289222 2294
rect 288986 -582 289222 -346
rect 288986 -902 289222 -666
rect 292686 689758 292922 689994
rect 292686 653758 292922 653994
rect 292686 617758 292922 617994
rect 292686 581758 292922 581994
rect 292686 545758 292922 545994
rect 292686 509758 292922 509994
rect 292686 473758 292922 473994
rect 292686 437758 292922 437994
rect 292686 401758 292922 401994
rect 292686 365758 292922 365994
rect 292686 329758 292922 329994
rect 292686 293758 292922 293994
rect 292686 257758 292922 257994
rect 292686 221758 292922 221994
rect 292686 185758 292922 185994
rect 292686 149758 292922 149994
rect 292686 113758 292922 113994
rect 292686 77758 292922 77994
rect 292686 41758 292922 41994
rect 292686 5758 292922 5994
rect 292686 -2502 292922 -2266
rect 292686 -2822 292922 -2586
rect 296386 693458 296622 693694
rect 296386 657458 296622 657694
rect 296386 621458 296622 621694
rect 296386 585458 296622 585694
rect 296386 549458 296622 549694
rect 296386 513458 296622 513694
rect 296386 477458 296622 477694
rect 296386 441458 296622 441694
rect 296386 405458 296622 405694
rect 296386 369458 296622 369694
rect 296386 333458 296622 333694
rect 296386 297458 296622 297694
rect 296386 261458 296622 261694
rect 296386 225458 296622 225694
rect 296386 189458 296622 189694
rect 296386 153458 296622 153694
rect 296386 117458 296622 117694
rect 296386 81458 296622 81694
rect 296386 45458 296622 45694
rect 296386 9458 296622 9694
rect 296386 -4422 296622 -4186
rect 296386 -4742 296622 -4506
rect 318086 711322 318322 711558
rect 318086 711002 318322 711238
rect 314386 709402 314622 709638
rect 314386 709082 314622 709318
rect 310686 707482 310922 707718
rect 310686 707162 310922 707398
rect 300086 697158 300322 697394
rect 300086 661158 300322 661394
rect 300086 625158 300322 625394
rect 300086 589158 300322 589394
rect 300086 553158 300322 553394
rect 300086 517158 300322 517394
rect 300086 481158 300322 481394
rect 300086 445158 300322 445394
rect 300086 409158 300322 409394
rect 300086 373158 300322 373394
rect 300086 337158 300322 337394
rect 300086 301158 300322 301394
rect 300086 265158 300322 265394
rect 300086 229158 300322 229394
rect 300086 193158 300322 193394
rect 300086 157158 300322 157394
rect 300086 121158 300322 121394
rect 300086 85158 300322 85394
rect 300086 49158 300322 49394
rect 300086 13158 300322 13394
rect 282086 -7302 282322 -7066
rect 282086 -7622 282322 -7386
rect 306986 705562 307222 705798
rect 306986 705242 307222 705478
rect 306986 668058 307222 668294
rect 306986 632058 307222 632294
rect 306986 596058 307222 596294
rect 306986 560058 307222 560294
rect 306986 524058 307222 524294
rect 306986 488058 307222 488294
rect 306986 452058 307222 452294
rect 306986 416058 307222 416294
rect 306986 380058 307222 380294
rect 306986 344058 307222 344294
rect 306986 308058 307222 308294
rect 306986 272058 307222 272294
rect 306986 236058 307222 236294
rect 306986 200058 307222 200294
rect 306986 164058 307222 164294
rect 306986 128058 307222 128294
rect 306986 92058 307222 92294
rect 306986 56058 307222 56294
rect 306986 20058 307222 20294
rect 306986 -1542 307222 -1306
rect 306986 -1862 307222 -1626
rect 310686 671758 310922 671994
rect 310686 635758 310922 635994
rect 310686 599758 310922 599994
rect 310686 563758 310922 563994
rect 310686 527758 310922 527994
rect 310686 491758 310922 491994
rect 310686 455758 310922 455994
rect 310686 419758 310922 419994
rect 310686 383758 310922 383994
rect 310686 347758 310922 347994
rect 310686 311758 310922 311994
rect 310686 275758 310922 275994
rect 310686 239758 310922 239994
rect 310686 203758 310922 203994
rect 310686 167758 310922 167994
rect 310686 131758 310922 131994
rect 310686 95758 310922 95994
rect 310686 59758 310922 59994
rect 310686 23758 310922 23994
rect 310686 -3462 310922 -3226
rect 310686 -3782 310922 -3546
rect 314386 675458 314622 675694
rect 314386 639458 314622 639694
rect 314386 603458 314622 603694
rect 314386 567458 314622 567694
rect 314386 531458 314622 531694
rect 314386 495458 314622 495694
rect 314386 459458 314622 459694
rect 314386 423458 314622 423694
rect 314386 387458 314622 387694
rect 314386 351458 314622 351694
rect 314386 315458 314622 315694
rect 314386 279458 314622 279694
rect 314386 243458 314622 243694
rect 314386 207458 314622 207694
rect 314386 171458 314622 171694
rect 314386 135458 314622 135694
rect 314386 99458 314622 99694
rect 314386 63458 314622 63694
rect 314386 27458 314622 27694
rect 314386 -5382 314622 -5146
rect 314386 -5702 314622 -5466
rect 336086 710362 336322 710598
rect 336086 710042 336322 710278
rect 332386 708442 332622 708678
rect 332386 708122 332622 708358
rect 328686 706522 328922 706758
rect 328686 706202 328922 706438
rect 318086 679158 318322 679394
rect 318086 643158 318322 643394
rect 318086 607158 318322 607394
rect 318086 571158 318322 571394
rect 318086 535158 318322 535394
rect 318086 499158 318322 499394
rect 318086 463158 318322 463394
rect 318086 427158 318322 427394
rect 318086 391158 318322 391394
rect 318086 355158 318322 355394
rect 318086 319158 318322 319394
rect 318086 283158 318322 283394
rect 318086 247158 318322 247394
rect 318086 211158 318322 211394
rect 318086 175158 318322 175394
rect 318086 139158 318322 139394
rect 318086 103158 318322 103394
rect 318086 67158 318322 67394
rect 318086 31158 318322 31394
rect 300086 -6342 300322 -6106
rect 300086 -6662 300322 -6426
rect 324986 704602 325222 704838
rect 324986 704282 325222 704518
rect 324986 686058 325222 686294
rect 324986 650058 325222 650294
rect 324986 614058 325222 614294
rect 324986 578058 325222 578294
rect 324986 542058 325222 542294
rect 324986 506058 325222 506294
rect 324986 470058 325222 470294
rect 324986 434058 325222 434294
rect 324986 398058 325222 398294
rect 324986 362058 325222 362294
rect 324986 326058 325222 326294
rect 324986 290058 325222 290294
rect 324986 254058 325222 254294
rect 324986 218058 325222 218294
rect 324986 182058 325222 182294
rect 324986 146058 325222 146294
rect 324986 110058 325222 110294
rect 324986 74058 325222 74294
rect 324986 38058 325222 38294
rect 324986 2058 325222 2294
rect 324986 -582 325222 -346
rect 324986 -902 325222 -666
rect 328686 689758 328922 689994
rect 328686 653758 328922 653994
rect 328686 617758 328922 617994
rect 328686 581758 328922 581994
rect 328686 545758 328922 545994
rect 328686 509758 328922 509994
rect 328686 473758 328922 473994
rect 328686 437758 328922 437994
rect 328686 401758 328922 401994
rect 328686 365758 328922 365994
rect 328686 329758 328922 329994
rect 328686 293758 328922 293994
rect 328686 257758 328922 257994
rect 328686 221758 328922 221994
rect 328686 185758 328922 185994
rect 328686 149758 328922 149994
rect 328686 113758 328922 113994
rect 328686 77758 328922 77994
rect 328686 41758 328922 41994
rect 328686 5758 328922 5994
rect 328686 -2502 328922 -2266
rect 328686 -2822 328922 -2586
rect 332386 693458 332622 693694
rect 332386 657458 332622 657694
rect 332386 621458 332622 621694
rect 332386 585458 332622 585694
rect 332386 549458 332622 549694
rect 332386 513458 332622 513694
rect 332386 477458 332622 477694
rect 332386 441458 332622 441694
rect 332386 405458 332622 405694
rect 332386 369458 332622 369694
rect 332386 333458 332622 333694
rect 332386 297458 332622 297694
rect 332386 261458 332622 261694
rect 332386 225458 332622 225694
rect 332386 189458 332622 189694
rect 332386 153458 332622 153694
rect 332386 117458 332622 117694
rect 332386 81458 332622 81694
rect 332386 45458 332622 45694
rect 332386 9458 332622 9694
rect 332386 -4422 332622 -4186
rect 332386 -4742 332622 -4506
rect 354086 711322 354322 711558
rect 354086 711002 354322 711238
rect 350386 709402 350622 709638
rect 350386 709082 350622 709318
rect 346686 707482 346922 707718
rect 346686 707162 346922 707398
rect 336086 697158 336322 697394
rect 336086 661158 336322 661394
rect 336086 625158 336322 625394
rect 336086 589158 336322 589394
rect 336086 553158 336322 553394
rect 336086 517158 336322 517394
rect 336086 481158 336322 481394
rect 336086 445158 336322 445394
rect 342986 705562 343222 705798
rect 342986 705242 343222 705478
rect 342986 668058 343222 668294
rect 342986 632058 343222 632294
rect 342986 596058 343222 596294
rect 342986 560058 343222 560294
rect 342986 524058 343222 524294
rect 342986 488058 343222 488294
rect 342986 452058 343222 452294
rect 346686 671758 346922 671994
rect 346686 635758 346922 635994
rect 346686 599758 346922 599994
rect 346686 563758 346922 563994
rect 346686 527758 346922 527994
rect 346686 491758 346922 491994
rect 346686 455758 346922 455994
rect 350386 675458 350622 675694
rect 350386 639458 350622 639694
rect 350386 603458 350622 603694
rect 350386 567458 350622 567694
rect 350386 531458 350622 531694
rect 350386 495458 350622 495694
rect 350386 459458 350622 459694
rect 372086 710362 372322 710598
rect 372086 710042 372322 710278
rect 368386 708442 368622 708678
rect 368386 708122 368622 708358
rect 364686 706522 364922 706758
rect 364686 706202 364922 706438
rect 354086 679158 354322 679394
rect 354086 643158 354322 643394
rect 354086 607158 354322 607394
rect 354086 571158 354322 571394
rect 354086 535158 354322 535394
rect 354086 499158 354322 499394
rect 354086 463158 354322 463394
rect 354086 427158 354322 427394
rect 360986 704602 361222 704838
rect 360986 704282 361222 704518
rect 360986 686058 361222 686294
rect 360986 650058 361222 650294
rect 360986 614058 361222 614294
rect 360986 578058 361222 578294
rect 360986 542058 361222 542294
rect 360986 506058 361222 506294
rect 360986 470058 361222 470294
rect 360986 434058 361222 434294
rect 364686 689758 364922 689994
rect 364686 653758 364922 653994
rect 364686 617758 364922 617994
rect 364686 581758 364922 581994
rect 364686 545758 364922 545994
rect 364686 509758 364922 509994
rect 364686 473758 364922 473994
rect 364686 437758 364922 437994
rect 368386 693458 368622 693694
rect 368386 657458 368622 657694
rect 368386 621458 368622 621694
rect 368386 585458 368622 585694
rect 368386 549458 368622 549694
rect 368386 513458 368622 513694
rect 368386 477458 368622 477694
rect 368386 441458 368622 441694
rect 390086 711322 390322 711558
rect 390086 711002 390322 711238
rect 386386 709402 386622 709638
rect 386386 709082 386622 709318
rect 382686 707482 382922 707718
rect 382686 707162 382922 707398
rect 372086 697158 372322 697394
rect 372086 661158 372322 661394
rect 372086 625158 372322 625394
rect 372086 589158 372322 589394
rect 372086 553158 372322 553394
rect 372086 517158 372322 517394
rect 372086 481158 372322 481394
rect 372086 445158 372322 445394
rect 378986 705562 379222 705798
rect 378986 705242 379222 705478
rect 378986 668058 379222 668294
rect 378986 632058 379222 632294
rect 378986 596058 379222 596294
rect 378986 560058 379222 560294
rect 378986 524058 379222 524294
rect 378986 488058 379222 488294
rect 378986 452058 379222 452294
rect 382686 671758 382922 671994
rect 382686 635758 382922 635994
rect 382686 599758 382922 599994
rect 382686 563758 382922 563994
rect 382686 527758 382922 527994
rect 382686 491758 382922 491994
rect 382686 455758 382922 455994
rect 386386 675458 386622 675694
rect 386386 639458 386622 639694
rect 386386 603458 386622 603694
rect 386386 567458 386622 567694
rect 386386 531458 386622 531694
rect 386386 495458 386622 495694
rect 386386 459458 386622 459694
rect 408086 710362 408322 710598
rect 408086 710042 408322 710278
rect 404386 708442 404622 708678
rect 404386 708122 404622 708358
rect 400686 706522 400922 706758
rect 400686 706202 400922 706438
rect 390086 679158 390322 679394
rect 390086 643158 390322 643394
rect 390086 607158 390322 607394
rect 390086 571158 390322 571394
rect 390086 535158 390322 535394
rect 390086 499158 390322 499394
rect 390086 463158 390322 463394
rect 390086 427158 390322 427394
rect 396986 704602 397222 704838
rect 396986 704282 397222 704518
rect 396986 686058 397222 686294
rect 396986 650058 397222 650294
rect 396986 614058 397222 614294
rect 396986 578058 397222 578294
rect 396986 542058 397222 542294
rect 396986 506058 397222 506294
rect 396986 470058 397222 470294
rect 396986 434058 397222 434294
rect 400686 689758 400922 689994
rect 400686 653758 400922 653994
rect 400686 617758 400922 617994
rect 400686 581758 400922 581994
rect 400686 545758 400922 545994
rect 400686 509758 400922 509994
rect 400686 473758 400922 473994
rect 400686 437758 400922 437994
rect 404386 693458 404622 693694
rect 404386 657458 404622 657694
rect 404386 621458 404622 621694
rect 404386 585458 404622 585694
rect 404386 549458 404622 549694
rect 404386 513458 404622 513694
rect 404386 477458 404622 477694
rect 404386 441458 404622 441694
rect 426086 711322 426322 711558
rect 426086 711002 426322 711238
rect 422386 709402 422622 709638
rect 422386 709082 422622 709318
rect 418686 707482 418922 707718
rect 418686 707162 418922 707398
rect 408086 697158 408322 697394
rect 408086 661158 408322 661394
rect 408086 625158 408322 625394
rect 408086 589158 408322 589394
rect 408086 553158 408322 553394
rect 408086 517158 408322 517394
rect 408086 481158 408322 481394
rect 408086 445158 408322 445394
rect 414986 705562 415222 705798
rect 414986 705242 415222 705478
rect 414986 668058 415222 668294
rect 414986 632058 415222 632294
rect 414986 596058 415222 596294
rect 414986 560058 415222 560294
rect 414986 524058 415222 524294
rect 414986 488058 415222 488294
rect 414986 452058 415222 452294
rect 418686 671758 418922 671994
rect 418686 635758 418922 635994
rect 418686 599758 418922 599994
rect 418686 563758 418922 563994
rect 418686 527758 418922 527994
rect 418686 491758 418922 491994
rect 418686 455758 418922 455994
rect 422386 675458 422622 675694
rect 422386 639458 422622 639694
rect 422386 603458 422622 603694
rect 422386 567458 422622 567694
rect 422386 531458 422622 531694
rect 422386 495458 422622 495694
rect 422386 459458 422622 459694
rect 444086 710362 444322 710598
rect 444086 710042 444322 710278
rect 440386 708442 440622 708678
rect 440386 708122 440622 708358
rect 436686 706522 436922 706758
rect 436686 706202 436922 706438
rect 426086 679158 426322 679394
rect 426086 643158 426322 643394
rect 426086 607158 426322 607394
rect 426086 571158 426322 571394
rect 426086 535158 426322 535394
rect 426086 499158 426322 499394
rect 426086 463158 426322 463394
rect 426086 427158 426322 427394
rect 432986 704602 433222 704838
rect 432986 704282 433222 704518
rect 432986 686058 433222 686294
rect 432986 650058 433222 650294
rect 432986 614058 433222 614294
rect 432986 578058 433222 578294
rect 432986 542058 433222 542294
rect 432986 506058 433222 506294
rect 432986 470058 433222 470294
rect 432986 434058 433222 434294
rect 436686 689758 436922 689994
rect 436686 653758 436922 653994
rect 436686 617758 436922 617994
rect 436686 581758 436922 581994
rect 436686 545758 436922 545994
rect 436686 509758 436922 509994
rect 436686 473758 436922 473994
rect 436686 437758 436922 437994
rect 440386 693458 440622 693694
rect 440386 657458 440622 657694
rect 440386 621458 440622 621694
rect 440386 585458 440622 585694
rect 440386 549458 440622 549694
rect 440386 513458 440622 513694
rect 440386 477458 440622 477694
rect 440386 441458 440622 441694
rect 462086 711322 462322 711558
rect 462086 711002 462322 711238
rect 458386 709402 458622 709638
rect 458386 709082 458622 709318
rect 454686 707482 454922 707718
rect 454686 707162 454922 707398
rect 444086 697158 444322 697394
rect 444086 661158 444322 661394
rect 444086 625158 444322 625394
rect 444086 589158 444322 589394
rect 444086 553158 444322 553394
rect 444086 517158 444322 517394
rect 444086 481158 444322 481394
rect 444086 445158 444322 445394
rect 450986 705562 451222 705798
rect 450986 705242 451222 705478
rect 450986 668058 451222 668294
rect 450986 632058 451222 632294
rect 450986 596058 451222 596294
rect 450986 560058 451222 560294
rect 450986 524058 451222 524294
rect 450986 488058 451222 488294
rect 450986 452058 451222 452294
rect 454686 671758 454922 671994
rect 454686 635758 454922 635994
rect 454686 599758 454922 599994
rect 454686 563758 454922 563994
rect 454686 527758 454922 527994
rect 454686 491758 454922 491994
rect 454686 455758 454922 455994
rect 458386 675458 458622 675694
rect 458386 639458 458622 639694
rect 458386 603458 458622 603694
rect 458386 567458 458622 567694
rect 458386 531458 458622 531694
rect 458386 495458 458622 495694
rect 458386 459458 458622 459694
rect 480086 710362 480322 710598
rect 480086 710042 480322 710278
rect 476386 708442 476622 708678
rect 476386 708122 476622 708358
rect 472686 706522 472922 706758
rect 472686 706202 472922 706438
rect 462086 679158 462322 679394
rect 462086 643158 462322 643394
rect 462086 607158 462322 607394
rect 462086 571158 462322 571394
rect 462086 535158 462322 535394
rect 462086 499158 462322 499394
rect 462086 463158 462322 463394
rect 462086 427158 462322 427394
rect 468986 704602 469222 704838
rect 468986 704282 469222 704518
rect 468986 686058 469222 686294
rect 468986 650058 469222 650294
rect 468986 614058 469222 614294
rect 468986 578058 469222 578294
rect 468986 542058 469222 542294
rect 468986 506058 469222 506294
rect 468986 470058 469222 470294
rect 468986 434058 469222 434294
rect 472686 689758 472922 689994
rect 472686 653758 472922 653994
rect 472686 617758 472922 617994
rect 472686 581758 472922 581994
rect 472686 545758 472922 545994
rect 472686 509758 472922 509994
rect 472686 473758 472922 473994
rect 472686 437758 472922 437994
rect 476386 693458 476622 693694
rect 476386 657458 476622 657694
rect 476386 621458 476622 621694
rect 476386 585458 476622 585694
rect 476386 549458 476622 549694
rect 476386 513458 476622 513694
rect 476386 477458 476622 477694
rect 476386 441458 476622 441694
rect 498086 711322 498322 711558
rect 498086 711002 498322 711238
rect 494386 709402 494622 709638
rect 494386 709082 494622 709318
rect 490686 707482 490922 707718
rect 490686 707162 490922 707398
rect 480086 697158 480322 697394
rect 480086 661158 480322 661394
rect 480086 625158 480322 625394
rect 480086 589158 480322 589394
rect 480086 553158 480322 553394
rect 480086 517158 480322 517394
rect 480086 481158 480322 481394
rect 480086 445158 480322 445394
rect 340328 416058 340564 416294
rect 476056 416058 476292 416294
rect 336086 409158 336322 409394
rect 480086 409158 480322 409394
rect 341008 398058 341244 398294
rect 475376 398058 475612 398294
rect 340328 380058 340564 380294
rect 476056 380058 476292 380294
rect 336086 373158 336322 373394
rect 480086 373158 480322 373394
rect 341008 362058 341244 362294
rect 475376 362058 475612 362294
rect 340328 344058 340564 344294
rect 476056 344058 476292 344294
rect 336086 337158 336322 337394
rect 336086 301158 336322 301394
rect 336086 265158 336322 265394
rect 336086 229158 336322 229394
rect 336086 193158 336322 193394
rect 336086 157158 336322 157394
rect 336086 121158 336322 121394
rect 336086 85158 336322 85394
rect 336086 49158 336322 49394
rect 336086 13158 336322 13394
rect 318086 -7302 318322 -7066
rect 318086 -7622 318322 -7386
rect 342986 308058 343222 308294
rect 342986 272058 343222 272294
rect 342986 236058 343222 236294
rect 342986 200058 343222 200294
rect 342986 164058 343222 164294
rect 342986 128058 343222 128294
rect 342986 92058 343222 92294
rect 342986 56058 343222 56294
rect 342986 20058 343222 20294
rect 342986 -1542 343222 -1306
rect 342986 -1862 343222 -1626
rect 346686 311758 346922 311994
rect 346686 275758 346922 275994
rect 346686 239758 346922 239994
rect 346686 203758 346922 203994
rect 346686 167758 346922 167994
rect 346686 131758 346922 131994
rect 346686 95758 346922 95994
rect 346686 59758 346922 59994
rect 346686 23758 346922 23994
rect 346686 -3462 346922 -3226
rect 346686 -3782 346922 -3546
rect 350386 315458 350622 315694
rect 350386 279458 350622 279694
rect 350386 243458 350622 243694
rect 350386 207458 350622 207694
rect 350386 171458 350622 171694
rect 350386 135458 350622 135694
rect 350386 99458 350622 99694
rect 350386 63458 350622 63694
rect 350386 27458 350622 27694
rect 350386 -5382 350622 -5146
rect 350386 -5702 350622 -5466
rect 354086 319158 354322 319394
rect 354086 283158 354322 283394
rect 354086 247158 354322 247394
rect 354086 211158 354322 211394
rect 354086 175158 354322 175394
rect 354086 139158 354322 139394
rect 354086 103158 354322 103394
rect 354086 67158 354322 67394
rect 354086 31158 354322 31394
rect 336086 -6342 336322 -6106
rect 336086 -6662 336322 -6426
rect 360986 326058 361222 326294
rect 360986 290058 361222 290294
rect 360986 254058 361222 254294
rect 360986 218058 361222 218294
rect 360986 182058 361222 182294
rect 360986 146058 361222 146294
rect 360986 110058 361222 110294
rect 360986 74058 361222 74294
rect 360986 38058 361222 38294
rect 360986 2058 361222 2294
rect 360986 -582 361222 -346
rect 360986 -902 361222 -666
rect 364686 329758 364922 329994
rect 364686 293758 364922 293994
rect 364686 257758 364922 257994
rect 364686 221758 364922 221994
rect 364686 185758 364922 185994
rect 364686 149758 364922 149994
rect 364686 113758 364922 113994
rect 364686 77758 364922 77994
rect 364686 41758 364922 41994
rect 364686 5758 364922 5994
rect 364686 -2502 364922 -2266
rect 364686 -2822 364922 -2586
rect 372086 337158 372322 337394
rect 368386 333458 368622 333694
rect 368386 297458 368622 297694
rect 368386 261458 368622 261694
rect 368386 225458 368622 225694
rect 368386 189458 368622 189694
rect 368386 153458 368622 153694
rect 368386 117458 368622 117694
rect 368386 81458 368622 81694
rect 368386 45458 368622 45694
rect 368386 9458 368622 9694
rect 368386 -4422 368622 -4186
rect 368386 -4742 368622 -4506
rect 372086 301158 372322 301394
rect 372086 265158 372322 265394
rect 372086 229158 372322 229394
rect 372086 193158 372322 193394
rect 372086 157158 372322 157394
rect 372086 121158 372322 121394
rect 372086 85158 372322 85394
rect 372086 49158 372322 49394
rect 372086 13158 372322 13394
rect 354086 -7302 354322 -7066
rect 354086 -7622 354322 -7386
rect 378986 308058 379222 308294
rect 378986 272058 379222 272294
rect 378986 236058 379222 236294
rect 378986 200058 379222 200294
rect 378986 164058 379222 164294
rect 378986 128058 379222 128294
rect 378986 92058 379222 92294
rect 378986 56058 379222 56294
rect 378986 20058 379222 20294
rect 378986 -1542 379222 -1306
rect 378986 -1862 379222 -1626
rect 382686 311758 382922 311994
rect 382686 275758 382922 275994
rect 382686 239758 382922 239994
rect 382686 203758 382922 203994
rect 382686 167758 382922 167994
rect 382686 131758 382922 131994
rect 382686 95758 382922 95994
rect 382686 59758 382922 59994
rect 382686 23758 382922 23994
rect 382686 -3462 382922 -3226
rect 382686 -3782 382922 -3546
rect 386386 315458 386622 315694
rect 386386 279458 386622 279694
rect 386386 243458 386622 243694
rect 386386 207458 386622 207694
rect 386386 171458 386622 171694
rect 386386 135458 386622 135694
rect 386386 99458 386622 99694
rect 386386 63458 386622 63694
rect 386386 27458 386622 27694
rect 386386 -5382 386622 -5146
rect 386386 -5702 386622 -5466
rect 390086 319158 390322 319394
rect 390086 283158 390322 283394
rect 390086 247158 390322 247394
rect 390086 211158 390322 211394
rect 390086 175158 390322 175394
rect 390086 139158 390322 139394
rect 390086 103158 390322 103394
rect 390086 67158 390322 67394
rect 390086 31158 390322 31394
rect 372086 -6342 372322 -6106
rect 372086 -6662 372322 -6426
rect 396986 326058 397222 326294
rect 396986 290058 397222 290294
rect 396986 254058 397222 254294
rect 396986 218058 397222 218294
rect 396986 182058 397222 182294
rect 396986 146058 397222 146294
rect 396986 110058 397222 110294
rect 396986 74058 397222 74294
rect 396986 38058 397222 38294
rect 396986 2058 397222 2294
rect 396986 -582 397222 -346
rect 396986 -902 397222 -666
rect 400686 329758 400922 329994
rect 400686 293758 400922 293994
rect 400686 257758 400922 257994
rect 400686 221758 400922 221994
rect 400686 185758 400922 185994
rect 400686 149758 400922 149994
rect 400686 113758 400922 113994
rect 400686 77758 400922 77994
rect 400686 41758 400922 41994
rect 400686 5758 400922 5994
rect 400686 -2502 400922 -2266
rect 400686 -2822 400922 -2586
rect 408086 337158 408322 337394
rect 404386 333458 404622 333694
rect 404386 297458 404622 297694
rect 404386 261458 404622 261694
rect 404386 225458 404622 225694
rect 404386 189458 404622 189694
rect 404386 153458 404622 153694
rect 404386 117458 404622 117694
rect 404386 81458 404622 81694
rect 404386 45458 404622 45694
rect 404386 9458 404622 9694
rect 404386 -4422 404622 -4186
rect 404386 -4742 404622 -4506
rect 408086 301158 408322 301394
rect 408086 265158 408322 265394
rect 408086 229158 408322 229394
rect 408086 193158 408322 193394
rect 408086 157158 408322 157394
rect 408086 121158 408322 121394
rect 408086 85158 408322 85394
rect 408086 49158 408322 49394
rect 408086 13158 408322 13394
rect 390086 -7302 390322 -7066
rect 390086 -7622 390322 -7386
rect 414986 308058 415222 308294
rect 414986 272058 415222 272294
rect 414986 236058 415222 236294
rect 414986 200058 415222 200294
rect 414986 164058 415222 164294
rect 414986 128058 415222 128294
rect 414986 92058 415222 92294
rect 414986 56058 415222 56294
rect 414986 20058 415222 20294
rect 414986 -1542 415222 -1306
rect 414986 -1862 415222 -1626
rect 418686 311758 418922 311994
rect 418686 275758 418922 275994
rect 418686 239758 418922 239994
rect 418686 203758 418922 203994
rect 418686 167758 418922 167994
rect 418686 131758 418922 131994
rect 418686 95758 418922 95994
rect 418686 59758 418922 59994
rect 418686 23758 418922 23994
rect 418686 -3462 418922 -3226
rect 418686 -3782 418922 -3546
rect 422386 315458 422622 315694
rect 422386 279458 422622 279694
rect 422386 243458 422622 243694
rect 422386 207458 422622 207694
rect 422386 171458 422622 171694
rect 422386 135458 422622 135694
rect 422386 99458 422622 99694
rect 422386 63458 422622 63694
rect 422386 27458 422622 27694
rect 422386 -5382 422622 -5146
rect 422386 -5702 422622 -5466
rect 426086 319158 426322 319394
rect 426086 283158 426322 283394
rect 426086 247158 426322 247394
rect 426086 211158 426322 211394
rect 426086 175158 426322 175394
rect 426086 139158 426322 139394
rect 426086 103158 426322 103394
rect 426086 67158 426322 67394
rect 426086 31158 426322 31394
rect 408086 -6342 408322 -6106
rect 408086 -6662 408322 -6426
rect 432986 326058 433222 326294
rect 432986 290058 433222 290294
rect 432986 254058 433222 254294
rect 432986 218058 433222 218294
rect 432986 182058 433222 182294
rect 432986 146058 433222 146294
rect 432986 110058 433222 110294
rect 432986 74058 433222 74294
rect 432986 38058 433222 38294
rect 432986 2058 433222 2294
rect 432986 -582 433222 -346
rect 432986 -902 433222 -666
rect 436686 329758 436922 329994
rect 436686 293758 436922 293994
rect 436686 257758 436922 257994
rect 436686 221758 436922 221994
rect 436686 185758 436922 185994
rect 436686 149758 436922 149994
rect 436686 113758 436922 113994
rect 436686 77758 436922 77994
rect 436686 41758 436922 41994
rect 436686 5758 436922 5994
rect 436686 -2502 436922 -2266
rect 436686 -2822 436922 -2586
rect 444086 337158 444322 337394
rect 440386 333458 440622 333694
rect 440386 297458 440622 297694
rect 440386 261458 440622 261694
rect 440386 225458 440622 225694
rect 440386 189458 440622 189694
rect 440386 153458 440622 153694
rect 440386 117458 440622 117694
rect 440386 81458 440622 81694
rect 440386 45458 440622 45694
rect 440386 9458 440622 9694
rect 440386 -4422 440622 -4186
rect 440386 -4742 440622 -4506
rect 444086 301158 444322 301394
rect 444086 265158 444322 265394
rect 444086 229158 444322 229394
rect 444086 193158 444322 193394
rect 444086 157158 444322 157394
rect 444086 121158 444322 121394
rect 444086 85158 444322 85394
rect 444086 49158 444322 49394
rect 444086 13158 444322 13394
rect 426086 -7302 426322 -7066
rect 426086 -7622 426322 -7386
rect 450986 308058 451222 308294
rect 450986 272058 451222 272294
rect 450986 236058 451222 236294
rect 450986 200058 451222 200294
rect 450986 164058 451222 164294
rect 450986 128058 451222 128294
rect 450986 92058 451222 92294
rect 450986 56058 451222 56294
rect 450986 20058 451222 20294
rect 450986 -1542 451222 -1306
rect 450986 -1862 451222 -1626
rect 454686 311758 454922 311994
rect 454686 275758 454922 275994
rect 454686 239758 454922 239994
rect 454686 203758 454922 203994
rect 454686 167758 454922 167994
rect 454686 131758 454922 131994
rect 454686 95758 454922 95994
rect 454686 59758 454922 59994
rect 454686 23758 454922 23994
rect 454686 -3462 454922 -3226
rect 454686 -3782 454922 -3546
rect 458386 315458 458622 315694
rect 458386 279458 458622 279694
rect 458386 243458 458622 243694
rect 458386 207458 458622 207694
rect 458386 171458 458622 171694
rect 458386 135458 458622 135694
rect 458386 99458 458622 99694
rect 458386 63458 458622 63694
rect 458386 27458 458622 27694
rect 458386 -5382 458622 -5146
rect 458386 -5702 458622 -5466
rect 462086 319158 462322 319394
rect 462086 283158 462322 283394
rect 462086 247158 462322 247394
rect 462086 211158 462322 211394
rect 462086 175158 462322 175394
rect 462086 139158 462322 139394
rect 462086 103158 462322 103394
rect 462086 67158 462322 67394
rect 462086 31158 462322 31394
rect 444086 -6342 444322 -6106
rect 444086 -6662 444322 -6426
rect 468986 326058 469222 326294
rect 468986 290058 469222 290294
rect 468986 254058 469222 254294
rect 468986 218058 469222 218294
rect 468986 182058 469222 182294
rect 468986 146058 469222 146294
rect 468986 110058 469222 110294
rect 468986 74058 469222 74294
rect 468986 38058 469222 38294
rect 468986 2058 469222 2294
rect 468986 -582 469222 -346
rect 468986 -902 469222 -666
rect 472686 329758 472922 329994
rect 472686 293758 472922 293994
rect 472686 257758 472922 257994
rect 472686 221758 472922 221994
rect 472686 185758 472922 185994
rect 472686 149758 472922 149994
rect 472686 113758 472922 113994
rect 472686 77758 472922 77994
rect 472686 41758 472922 41994
rect 472686 5758 472922 5994
rect 472686 -2502 472922 -2266
rect 472686 -2822 472922 -2586
rect 476386 333458 476622 333694
rect 476386 297458 476622 297694
rect 476386 261458 476622 261694
rect 476386 225458 476622 225694
rect 476386 189458 476622 189694
rect 476386 153458 476622 153694
rect 476386 117458 476622 117694
rect 476386 81458 476622 81694
rect 476386 45458 476622 45694
rect 476386 9458 476622 9694
rect 476386 -4422 476622 -4186
rect 476386 -4742 476622 -4506
rect 480086 337158 480322 337394
rect 480086 301158 480322 301394
rect 480086 265158 480322 265394
rect 480086 229158 480322 229394
rect 480086 193158 480322 193394
rect 480086 157158 480322 157394
rect 480086 121158 480322 121394
rect 480086 85158 480322 85394
rect 480086 49158 480322 49394
rect 480086 13158 480322 13394
rect 462086 -7302 462322 -7066
rect 462086 -7622 462322 -7386
rect 486986 705562 487222 705798
rect 486986 705242 487222 705478
rect 486986 668058 487222 668294
rect 486986 632058 487222 632294
rect 486986 596058 487222 596294
rect 486986 560058 487222 560294
rect 486986 524058 487222 524294
rect 486986 488058 487222 488294
rect 486986 452058 487222 452294
rect 486986 416058 487222 416294
rect 486986 380058 487222 380294
rect 486986 344058 487222 344294
rect 486986 308058 487222 308294
rect 486986 272058 487222 272294
rect 486986 236058 487222 236294
rect 486986 200058 487222 200294
rect 486986 164058 487222 164294
rect 486986 128058 487222 128294
rect 486986 92058 487222 92294
rect 486986 56058 487222 56294
rect 486986 20058 487222 20294
rect 486986 -1542 487222 -1306
rect 486986 -1862 487222 -1626
rect 490686 671758 490922 671994
rect 490686 635758 490922 635994
rect 490686 599758 490922 599994
rect 490686 563758 490922 563994
rect 490686 527758 490922 527994
rect 490686 491758 490922 491994
rect 490686 455758 490922 455994
rect 490686 419758 490922 419994
rect 490686 383758 490922 383994
rect 490686 347758 490922 347994
rect 490686 311758 490922 311994
rect 490686 275758 490922 275994
rect 490686 239758 490922 239994
rect 490686 203758 490922 203994
rect 490686 167758 490922 167994
rect 490686 131758 490922 131994
rect 490686 95758 490922 95994
rect 490686 59758 490922 59994
rect 490686 23758 490922 23994
rect 490686 -3462 490922 -3226
rect 490686 -3782 490922 -3546
rect 494386 675458 494622 675694
rect 494386 639458 494622 639694
rect 494386 603458 494622 603694
rect 494386 567458 494622 567694
rect 494386 531458 494622 531694
rect 494386 495458 494622 495694
rect 494386 459458 494622 459694
rect 494386 423458 494622 423694
rect 494386 387458 494622 387694
rect 494386 351458 494622 351694
rect 494386 315458 494622 315694
rect 494386 279458 494622 279694
rect 494386 243458 494622 243694
rect 494386 207458 494622 207694
rect 494386 171458 494622 171694
rect 494386 135458 494622 135694
rect 494386 99458 494622 99694
rect 494386 63458 494622 63694
rect 494386 27458 494622 27694
rect 494386 -5382 494622 -5146
rect 494386 -5702 494622 -5466
rect 516086 710362 516322 710598
rect 516086 710042 516322 710278
rect 512386 708442 512622 708678
rect 512386 708122 512622 708358
rect 508686 706522 508922 706758
rect 508686 706202 508922 706438
rect 498086 679158 498322 679394
rect 498086 643158 498322 643394
rect 498086 607158 498322 607394
rect 498086 571158 498322 571394
rect 498086 535158 498322 535394
rect 498086 499158 498322 499394
rect 498086 463158 498322 463394
rect 498086 427158 498322 427394
rect 498086 391158 498322 391394
rect 498086 355158 498322 355394
rect 498086 319158 498322 319394
rect 498086 283158 498322 283394
rect 498086 247158 498322 247394
rect 498086 211158 498322 211394
rect 498086 175158 498322 175394
rect 498086 139158 498322 139394
rect 498086 103158 498322 103394
rect 498086 67158 498322 67394
rect 498086 31158 498322 31394
rect 480086 -6342 480322 -6106
rect 480086 -6662 480322 -6426
rect 504986 704602 505222 704838
rect 504986 704282 505222 704518
rect 504986 686058 505222 686294
rect 504986 650058 505222 650294
rect 504986 614058 505222 614294
rect 504986 578058 505222 578294
rect 504986 542058 505222 542294
rect 504986 506058 505222 506294
rect 504986 470058 505222 470294
rect 504986 434058 505222 434294
rect 504986 398058 505222 398294
rect 504986 362058 505222 362294
rect 504986 326058 505222 326294
rect 504986 290058 505222 290294
rect 504986 254058 505222 254294
rect 504986 218058 505222 218294
rect 504986 182058 505222 182294
rect 504986 146058 505222 146294
rect 504986 110058 505222 110294
rect 504986 74058 505222 74294
rect 504986 38058 505222 38294
rect 504986 2058 505222 2294
rect 504986 -582 505222 -346
rect 504986 -902 505222 -666
rect 508686 689758 508922 689994
rect 508686 653758 508922 653994
rect 508686 617758 508922 617994
rect 508686 581758 508922 581994
rect 508686 545758 508922 545994
rect 508686 509758 508922 509994
rect 508686 473758 508922 473994
rect 508686 437758 508922 437994
rect 508686 401758 508922 401994
rect 508686 365758 508922 365994
rect 508686 329758 508922 329994
rect 508686 293758 508922 293994
rect 508686 257758 508922 257994
rect 508686 221758 508922 221994
rect 508686 185758 508922 185994
rect 508686 149758 508922 149994
rect 508686 113758 508922 113994
rect 508686 77758 508922 77994
rect 508686 41758 508922 41994
rect 508686 5758 508922 5994
rect 508686 -2502 508922 -2266
rect 508686 -2822 508922 -2586
rect 512386 693458 512622 693694
rect 512386 657458 512622 657694
rect 512386 621458 512622 621694
rect 512386 585458 512622 585694
rect 512386 549458 512622 549694
rect 512386 513458 512622 513694
rect 512386 477458 512622 477694
rect 512386 441458 512622 441694
rect 512386 405458 512622 405694
rect 512386 369458 512622 369694
rect 512386 333458 512622 333694
rect 512386 297458 512622 297694
rect 512386 261458 512622 261694
rect 512386 225458 512622 225694
rect 512386 189458 512622 189694
rect 512386 153458 512622 153694
rect 512386 117458 512622 117694
rect 512386 81458 512622 81694
rect 512386 45458 512622 45694
rect 512386 9458 512622 9694
rect 512386 -4422 512622 -4186
rect 512386 -4742 512622 -4506
rect 534086 711322 534322 711558
rect 534086 711002 534322 711238
rect 530386 709402 530622 709638
rect 530386 709082 530622 709318
rect 526686 707482 526922 707718
rect 526686 707162 526922 707398
rect 516086 697158 516322 697394
rect 516086 661158 516322 661394
rect 516086 625158 516322 625394
rect 516086 589158 516322 589394
rect 516086 553158 516322 553394
rect 516086 517158 516322 517394
rect 516086 481158 516322 481394
rect 516086 445158 516322 445394
rect 516086 409158 516322 409394
rect 516086 373158 516322 373394
rect 516086 337158 516322 337394
rect 516086 301158 516322 301394
rect 516086 265158 516322 265394
rect 516086 229158 516322 229394
rect 516086 193158 516322 193394
rect 516086 157158 516322 157394
rect 516086 121158 516322 121394
rect 516086 85158 516322 85394
rect 516086 49158 516322 49394
rect 516086 13158 516322 13394
rect 498086 -7302 498322 -7066
rect 498086 -7622 498322 -7386
rect 522986 705562 523222 705798
rect 522986 705242 523222 705478
rect 522986 668058 523222 668294
rect 522986 632058 523222 632294
rect 522986 596058 523222 596294
rect 522986 560058 523222 560294
rect 522986 524058 523222 524294
rect 522986 488058 523222 488294
rect 522986 452058 523222 452294
rect 522986 416058 523222 416294
rect 522986 380058 523222 380294
rect 522986 344058 523222 344294
rect 522986 308058 523222 308294
rect 522986 272058 523222 272294
rect 522986 236058 523222 236294
rect 522986 200058 523222 200294
rect 522986 164058 523222 164294
rect 522986 128058 523222 128294
rect 522986 92058 523222 92294
rect 522986 56058 523222 56294
rect 522986 20058 523222 20294
rect 522986 -1542 523222 -1306
rect 522986 -1862 523222 -1626
rect 526686 671758 526922 671994
rect 526686 635758 526922 635994
rect 526686 599758 526922 599994
rect 526686 563758 526922 563994
rect 526686 527758 526922 527994
rect 526686 491758 526922 491994
rect 526686 455758 526922 455994
rect 526686 419758 526922 419994
rect 526686 383758 526922 383994
rect 526686 347758 526922 347994
rect 526686 311758 526922 311994
rect 526686 275758 526922 275994
rect 526686 239758 526922 239994
rect 526686 203758 526922 203994
rect 526686 167758 526922 167994
rect 526686 131758 526922 131994
rect 526686 95758 526922 95994
rect 526686 59758 526922 59994
rect 526686 23758 526922 23994
rect 526686 -3462 526922 -3226
rect 526686 -3782 526922 -3546
rect 530386 675458 530622 675694
rect 530386 639458 530622 639694
rect 530386 603458 530622 603694
rect 530386 567458 530622 567694
rect 530386 531458 530622 531694
rect 530386 495458 530622 495694
rect 530386 459458 530622 459694
rect 530386 423458 530622 423694
rect 530386 387458 530622 387694
rect 530386 351458 530622 351694
rect 530386 315458 530622 315694
rect 530386 279458 530622 279694
rect 530386 243458 530622 243694
rect 530386 207458 530622 207694
rect 530386 171458 530622 171694
rect 530386 135458 530622 135694
rect 530386 99458 530622 99694
rect 530386 63458 530622 63694
rect 530386 27458 530622 27694
rect 530386 -5382 530622 -5146
rect 530386 -5702 530622 -5466
rect 552086 710362 552322 710598
rect 552086 710042 552322 710278
rect 548386 708442 548622 708678
rect 548386 708122 548622 708358
rect 544686 706522 544922 706758
rect 544686 706202 544922 706438
rect 534086 679158 534322 679394
rect 534086 643158 534322 643394
rect 534086 607158 534322 607394
rect 534086 571158 534322 571394
rect 534086 535158 534322 535394
rect 534086 499158 534322 499394
rect 534086 463158 534322 463394
rect 534086 427158 534322 427394
rect 534086 391158 534322 391394
rect 534086 355158 534322 355394
rect 534086 319158 534322 319394
rect 534086 283158 534322 283394
rect 534086 247158 534322 247394
rect 534086 211158 534322 211394
rect 534086 175158 534322 175394
rect 534086 139158 534322 139394
rect 534086 103158 534322 103394
rect 534086 67158 534322 67394
rect 534086 31158 534322 31394
rect 516086 -6342 516322 -6106
rect 516086 -6662 516322 -6426
rect 540986 704602 541222 704838
rect 540986 704282 541222 704518
rect 540986 686058 541222 686294
rect 540986 650058 541222 650294
rect 540986 614058 541222 614294
rect 540986 578058 541222 578294
rect 540986 542058 541222 542294
rect 540986 506058 541222 506294
rect 540986 470058 541222 470294
rect 540986 434058 541222 434294
rect 540986 398058 541222 398294
rect 540986 362058 541222 362294
rect 540986 326058 541222 326294
rect 540986 290058 541222 290294
rect 540986 254058 541222 254294
rect 540986 218058 541222 218294
rect 540986 182058 541222 182294
rect 540986 146058 541222 146294
rect 540986 110058 541222 110294
rect 540986 74058 541222 74294
rect 540986 38058 541222 38294
rect 540986 2058 541222 2294
rect 540986 -582 541222 -346
rect 540986 -902 541222 -666
rect 544686 689758 544922 689994
rect 544686 653758 544922 653994
rect 544686 617758 544922 617994
rect 544686 581758 544922 581994
rect 544686 545758 544922 545994
rect 544686 509758 544922 509994
rect 544686 473758 544922 473994
rect 544686 437758 544922 437994
rect 544686 401758 544922 401994
rect 544686 365758 544922 365994
rect 544686 329758 544922 329994
rect 544686 293758 544922 293994
rect 544686 257758 544922 257994
rect 544686 221758 544922 221994
rect 544686 185758 544922 185994
rect 544686 149758 544922 149994
rect 544686 113758 544922 113994
rect 544686 77758 544922 77994
rect 544686 41758 544922 41994
rect 544686 5758 544922 5994
rect 544686 -2502 544922 -2266
rect 544686 -2822 544922 -2586
rect 548386 693458 548622 693694
rect 548386 657458 548622 657694
rect 548386 621458 548622 621694
rect 548386 585458 548622 585694
rect 548386 549458 548622 549694
rect 548386 513458 548622 513694
rect 548386 477458 548622 477694
rect 548386 441458 548622 441694
rect 548386 405458 548622 405694
rect 548386 369458 548622 369694
rect 548386 333458 548622 333694
rect 548386 297458 548622 297694
rect 548386 261458 548622 261694
rect 548386 225458 548622 225694
rect 548386 189458 548622 189694
rect 548386 153458 548622 153694
rect 548386 117458 548622 117694
rect 548386 81458 548622 81694
rect 548386 45458 548622 45694
rect 548386 9458 548622 9694
rect 548386 -4422 548622 -4186
rect 548386 -4742 548622 -4506
rect 570086 711322 570322 711558
rect 570086 711002 570322 711238
rect 566386 709402 566622 709638
rect 566386 709082 566622 709318
rect 562686 707482 562922 707718
rect 562686 707162 562922 707398
rect 552086 697158 552322 697394
rect 552086 661158 552322 661394
rect 552086 625158 552322 625394
rect 552086 589158 552322 589394
rect 552086 553158 552322 553394
rect 552086 517158 552322 517394
rect 552086 481158 552322 481394
rect 552086 445158 552322 445394
rect 552086 409158 552322 409394
rect 552086 373158 552322 373394
rect 552086 337158 552322 337394
rect 552086 301158 552322 301394
rect 552086 265158 552322 265394
rect 552086 229158 552322 229394
rect 552086 193158 552322 193394
rect 552086 157158 552322 157394
rect 552086 121158 552322 121394
rect 552086 85158 552322 85394
rect 552086 49158 552322 49394
rect 552086 13158 552322 13394
rect 534086 -7302 534322 -7066
rect 534086 -7622 534322 -7386
rect 558986 705562 559222 705798
rect 558986 705242 559222 705478
rect 558986 668058 559222 668294
rect 558986 632058 559222 632294
rect 558986 596058 559222 596294
rect 558986 560058 559222 560294
rect 558986 524058 559222 524294
rect 558986 488058 559222 488294
rect 558986 452058 559222 452294
rect 558986 416058 559222 416294
rect 558986 380058 559222 380294
rect 558986 344058 559222 344294
rect 558986 308058 559222 308294
rect 558986 272058 559222 272294
rect 558986 236058 559222 236294
rect 558986 200058 559222 200294
rect 558986 164058 559222 164294
rect 558986 128058 559222 128294
rect 558986 92058 559222 92294
rect 558986 56058 559222 56294
rect 558986 20058 559222 20294
rect 558986 -1542 559222 -1306
rect 558986 -1862 559222 -1626
rect 562686 671758 562922 671994
rect 562686 635758 562922 635994
rect 562686 599758 562922 599994
rect 562686 563758 562922 563994
rect 562686 527758 562922 527994
rect 562686 491758 562922 491994
rect 562686 455758 562922 455994
rect 562686 419758 562922 419994
rect 562686 383758 562922 383994
rect 562686 347758 562922 347994
rect 562686 311758 562922 311994
rect 562686 275758 562922 275994
rect 562686 239758 562922 239994
rect 562686 203758 562922 203994
rect 562686 167758 562922 167994
rect 562686 131758 562922 131994
rect 562686 95758 562922 95994
rect 562686 59758 562922 59994
rect 562686 23758 562922 23994
rect 562686 -3462 562922 -3226
rect 562686 -3782 562922 -3546
rect 566386 675458 566622 675694
rect 566386 639458 566622 639694
rect 566386 603458 566622 603694
rect 566386 567458 566622 567694
rect 566386 531458 566622 531694
rect 566386 495458 566622 495694
rect 566386 459458 566622 459694
rect 566386 423458 566622 423694
rect 566386 387458 566622 387694
rect 566386 351458 566622 351694
rect 566386 315458 566622 315694
rect 566386 279458 566622 279694
rect 566386 243458 566622 243694
rect 566386 207458 566622 207694
rect 566386 171458 566622 171694
rect 566386 135458 566622 135694
rect 566386 99458 566622 99694
rect 566386 63458 566622 63694
rect 566386 27458 566622 27694
rect 566386 -5382 566622 -5146
rect 566386 -5702 566622 -5466
rect 592062 711322 592298 711558
rect 592382 711322 592618 711558
rect 592062 711002 592298 711238
rect 592382 711002 592618 711238
rect 591102 710362 591338 710598
rect 591422 710362 591658 710598
rect 591102 710042 591338 710278
rect 591422 710042 591658 710278
rect 590142 709402 590378 709638
rect 590462 709402 590698 709638
rect 590142 709082 590378 709318
rect 590462 709082 590698 709318
rect 589182 708442 589418 708678
rect 589502 708442 589738 708678
rect 589182 708122 589418 708358
rect 589502 708122 589738 708358
rect 588222 707482 588458 707718
rect 588542 707482 588778 707718
rect 588222 707162 588458 707398
rect 588542 707162 588778 707398
rect 580686 706522 580922 706758
rect 580686 706202 580922 706438
rect 570086 679158 570322 679394
rect 570086 643158 570322 643394
rect 570086 607158 570322 607394
rect 570086 571158 570322 571394
rect 570086 535158 570322 535394
rect 570086 499158 570322 499394
rect 570086 463158 570322 463394
rect 570086 427158 570322 427394
rect 570086 391158 570322 391394
rect 570086 355158 570322 355394
rect 570086 319158 570322 319394
rect 570086 283158 570322 283394
rect 570086 247158 570322 247394
rect 570086 211158 570322 211394
rect 570086 175158 570322 175394
rect 570086 139158 570322 139394
rect 570086 103158 570322 103394
rect 570086 67158 570322 67394
rect 570086 31158 570322 31394
rect 552086 -6342 552322 -6106
rect 552086 -6662 552322 -6426
rect 576986 704602 577222 704838
rect 576986 704282 577222 704518
rect 576986 686058 577222 686294
rect 576986 650058 577222 650294
rect 576986 614058 577222 614294
rect 576986 578058 577222 578294
rect 576986 542058 577222 542294
rect 576986 506058 577222 506294
rect 576986 470058 577222 470294
rect 576986 434058 577222 434294
rect 576986 398058 577222 398294
rect 576986 362058 577222 362294
rect 576986 326058 577222 326294
rect 576986 290058 577222 290294
rect 576986 254058 577222 254294
rect 576986 218058 577222 218294
rect 576986 182058 577222 182294
rect 576986 146058 577222 146294
rect 576986 110058 577222 110294
rect 576986 74058 577222 74294
rect 576986 38058 577222 38294
rect 576986 2058 577222 2294
rect 576986 -582 577222 -346
rect 576986 -902 577222 -666
rect 587262 706522 587498 706758
rect 587582 706522 587818 706758
rect 587262 706202 587498 706438
rect 587582 706202 587818 706438
rect 586302 705562 586538 705798
rect 586622 705562 586858 705798
rect 586302 705242 586538 705478
rect 586622 705242 586858 705478
rect 580686 689758 580922 689994
rect 580686 653758 580922 653994
rect 580686 617758 580922 617994
rect 580686 581758 580922 581994
rect 580686 545758 580922 545994
rect 580686 509758 580922 509994
rect 580686 473758 580922 473994
rect 580686 437758 580922 437994
rect 580686 401758 580922 401994
rect 580686 365758 580922 365994
rect 580686 329758 580922 329994
rect 580686 293758 580922 293994
rect 580686 257758 580922 257994
rect 580686 221758 580922 221994
rect 580686 185758 580922 185994
rect 580686 149758 580922 149994
rect 580686 113758 580922 113994
rect 580686 77758 580922 77994
rect 580686 41758 580922 41994
rect 580686 5758 580922 5994
rect 585342 704602 585578 704838
rect 585662 704602 585898 704838
rect 585342 704282 585578 704518
rect 585662 704282 585898 704518
rect 585342 686058 585578 686294
rect 585662 686058 585898 686294
rect 585342 650058 585578 650294
rect 585662 650058 585898 650294
rect 585342 614058 585578 614294
rect 585662 614058 585898 614294
rect 585342 578058 585578 578294
rect 585662 578058 585898 578294
rect 585342 542058 585578 542294
rect 585662 542058 585898 542294
rect 585342 506058 585578 506294
rect 585662 506058 585898 506294
rect 585342 470058 585578 470294
rect 585662 470058 585898 470294
rect 585342 434058 585578 434294
rect 585662 434058 585898 434294
rect 585342 398058 585578 398294
rect 585662 398058 585898 398294
rect 585342 362058 585578 362294
rect 585662 362058 585898 362294
rect 585342 326058 585578 326294
rect 585662 326058 585898 326294
rect 585342 290058 585578 290294
rect 585662 290058 585898 290294
rect 585342 254058 585578 254294
rect 585662 254058 585898 254294
rect 585342 218058 585578 218294
rect 585662 218058 585898 218294
rect 585342 182058 585578 182294
rect 585662 182058 585898 182294
rect 585342 146058 585578 146294
rect 585662 146058 585898 146294
rect 585342 110058 585578 110294
rect 585662 110058 585898 110294
rect 585342 74058 585578 74294
rect 585662 74058 585898 74294
rect 585342 38058 585578 38294
rect 585662 38058 585898 38294
rect 585342 2058 585578 2294
rect 585662 2058 585898 2294
rect 585342 -582 585578 -346
rect 585662 -582 585898 -346
rect 585342 -902 585578 -666
rect 585662 -902 585898 -666
rect 586302 668058 586538 668294
rect 586622 668058 586858 668294
rect 586302 632058 586538 632294
rect 586622 632058 586858 632294
rect 586302 596058 586538 596294
rect 586622 596058 586858 596294
rect 586302 560058 586538 560294
rect 586622 560058 586858 560294
rect 586302 524058 586538 524294
rect 586622 524058 586858 524294
rect 586302 488058 586538 488294
rect 586622 488058 586858 488294
rect 586302 452058 586538 452294
rect 586622 452058 586858 452294
rect 586302 416058 586538 416294
rect 586622 416058 586858 416294
rect 586302 380058 586538 380294
rect 586622 380058 586858 380294
rect 586302 344058 586538 344294
rect 586622 344058 586858 344294
rect 586302 308058 586538 308294
rect 586622 308058 586858 308294
rect 586302 272058 586538 272294
rect 586622 272058 586858 272294
rect 586302 236058 586538 236294
rect 586622 236058 586858 236294
rect 586302 200058 586538 200294
rect 586622 200058 586858 200294
rect 586302 164058 586538 164294
rect 586622 164058 586858 164294
rect 586302 128058 586538 128294
rect 586622 128058 586858 128294
rect 586302 92058 586538 92294
rect 586622 92058 586858 92294
rect 586302 56058 586538 56294
rect 586622 56058 586858 56294
rect 586302 20058 586538 20294
rect 586622 20058 586858 20294
rect 586302 -1542 586538 -1306
rect 586622 -1542 586858 -1306
rect 586302 -1862 586538 -1626
rect 586622 -1862 586858 -1626
rect 587262 689758 587498 689994
rect 587582 689758 587818 689994
rect 587262 653758 587498 653994
rect 587582 653758 587818 653994
rect 587262 617758 587498 617994
rect 587582 617758 587818 617994
rect 587262 581758 587498 581994
rect 587582 581758 587818 581994
rect 587262 545758 587498 545994
rect 587582 545758 587818 545994
rect 587262 509758 587498 509994
rect 587582 509758 587818 509994
rect 587262 473758 587498 473994
rect 587582 473758 587818 473994
rect 587262 437758 587498 437994
rect 587582 437758 587818 437994
rect 587262 401758 587498 401994
rect 587582 401758 587818 401994
rect 587262 365758 587498 365994
rect 587582 365758 587818 365994
rect 587262 329758 587498 329994
rect 587582 329758 587818 329994
rect 587262 293758 587498 293994
rect 587582 293758 587818 293994
rect 587262 257758 587498 257994
rect 587582 257758 587818 257994
rect 587262 221758 587498 221994
rect 587582 221758 587818 221994
rect 587262 185758 587498 185994
rect 587582 185758 587818 185994
rect 587262 149758 587498 149994
rect 587582 149758 587818 149994
rect 587262 113758 587498 113994
rect 587582 113758 587818 113994
rect 587262 77758 587498 77994
rect 587582 77758 587818 77994
rect 587262 41758 587498 41994
rect 587582 41758 587818 41994
rect 587262 5758 587498 5994
rect 587582 5758 587818 5994
rect 580686 -2502 580922 -2266
rect 580686 -2822 580922 -2586
rect 587262 -2502 587498 -2266
rect 587582 -2502 587818 -2266
rect 587262 -2822 587498 -2586
rect 587582 -2822 587818 -2586
rect 588222 671758 588458 671994
rect 588542 671758 588778 671994
rect 588222 635758 588458 635994
rect 588542 635758 588778 635994
rect 588222 599758 588458 599994
rect 588542 599758 588778 599994
rect 588222 563758 588458 563994
rect 588542 563758 588778 563994
rect 588222 527758 588458 527994
rect 588542 527758 588778 527994
rect 588222 491758 588458 491994
rect 588542 491758 588778 491994
rect 588222 455758 588458 455994
rect 588542 455758 588778 455994
rect 588222 419758 588458 419994
rect 588542 419758 588778 419994
rect 588222 383758 588458 383994
rect 588542 383758 588778 383994
rect 588222 347758 588458 347994
rect 588542 347758 588778 347994
rect 588222 311758 588458 311994
rect 588542 311758 588778 311994
rect 588222 275758 588458 275994
rect 588542 275758 588778 275994
rect 588222 239758 588458 239994
rect 588542 239758 588778 239994
rect 588222 203758 588458 203994
rect 588542 203758 588778 203994
rect 588222 167758 588458 167994
rect 588542 167758 588778 167994
rect 588222 131758 588458 131994
rect 588542 131758 588778 131994
rect 588222 95758 588458 95994
rect 588542 95758 588778 95994
rect 588222 59758 588458 59994
rect 588542 59758 588778 59994
rect 588222 23758 588458 23994
rect 588542 23758 588778 23994
rect 588222 -3462 588458 -3226
rect 588542 -3462 588778 -3226
rect 588222 -3782 588458 -3546
rect 588542 -3782 588778 -3546
rect 589182 693458 589418 693694
rect 589502 693458 589738 693694
rect 589182 657458 589418 657694
rect 589502 657458 589738 657694
rect 589182 621458 589418 621694
rect 589502 621458 589738 621694
rect 589182 585458 589418 585694
rect 589502 585458 589738 585694
rect 589182 549458 589418 549694
rect 589502 549458 589738 549694
rect 589182 513458 589418 513694
rect 589502 513458 589738 513694
rect 589182 477458 589418 477694
rect 589502 477458 589738 477694
rect 589182 441458 589418 441694
rect 589502 441458 589738 441694
rect 589182 405458 589418 405694
rect 589502 405458 589738 405694
rect 589182 369458 589418 369694
rect 589502 369458 589738 369694
rect 589182 333458 589418 333694
rect 589502 333458 589738 333694
rect 589182 297458 589418 297694
rect 589502 297458 589738 297694
rect 589182 261458 589418 261694
rect 589502 261458 589738 261694
rect 589182 225458 589418 225694
rect 589502 225458 589738 225694
rect 589182 189458 589418 189694
rect 589502 189458 589738 189694
rect 589182 153458 589418 153694
rect 589502 153458 589738 153694
rect 589182 117458 589418 117694
rect 589502 117458 589738 117694
rect 589182 81458 589418 81694
rect 589502 81458 589738 81694
rect 589182 45458 589418 45694
rect 589502 45458 589738 45694
rect 589182 9458 589418 9694
rect 589502 9458 589738 9694
rect 589182 -4422 589418 -4186
rect 589502 -4422 589738 -4186
rect 589182 -4742 589418 -4506
rect 589502 -4742 589738 -4506
rect 590142 675458 590378 675694
rect 590462 675458 590698 675694
rect 590142 639458 590378 639694
rect 590462 639458 590698 639694
rect 590142 603458 590378 603694
rect 590462 603458 590698 603694
rect 590142 567458 590378 567694
rect 590462 567458 590698 567694
rect 590142 531458 590378 531694
rect 590462 531458 590698 531694
rect 590142 495458 590378 495694
rect 590462 495458 590698 495694
rect 590142 459458 590378 459694
rect 590462 459458 590698 459694
rect 590142 423458 590378 423694
rect 590462 423458 590698 423694
rect 590142 387458 590378 387694
rect 590462 387458 590698 387694
rect 590142 351458 590378 351694
rect 590462 351458 590698 351694
rect 590142 315458 590378 315694
rect 590462 315458 590698 315694
rect 590142 279458 590378 279694
rect 590462 279458 590698 279694
rect 590142 243458 590378 243694
rect 590462 243458 590698 243694
rect 590142 207458 590378 207694
rect 590462 207458 590698 207694
rect 590142 171458 590378 171694
rect 590462 171458 590698 171694
rect 590142 135458 590378 135694
rect 590462 135458 590698 135694
rect 590142 99458 590378 99694
rect 590462 99458 590698 99694
rect 590142 63458 590378 63694
rect 590462 63458 590698 63694
rect 590142 27458 590378 27694
rect 590462 27458 590698 27694
rect 590142 -5382 590378 -5146
rect 590462 -5382 590698 -5146
rect 590142 -5702 590378 -5466
rect 590462 -5702 590698 -5466
rect 591102 697158 591338 697394
rect 591422 697158 591658 697394
rect 591102 661158 591338 661394
rect 591422 661158 591658 661394
rect 591102 625158 591338 625394
rect 591422 625158 591658 625394
rect 591102 589158 591338 589394
rect 591422 589158 591658 589394
rect 591102 553158 591338 553394
rect 591422 553158 591658 553394
rect 591102 517158 591338 517394
rect 591422 517158 591658 517394
rect 591102 481158 591338 481394
rect 591422 481158 591658 481394
rect 591102 445158 591338 445394
rect 591422 445158 591658 445394
rect 591102 409158 591338 409394
rect 591422 409158 591658 409394
rect 591102 373158 591338 373394
rect 591422 373158 591658 373394
rect 591102 337158 591338 337394
rect 591422 337158 591658 337394
rect 591102 301158 591338 301394
rect 591422 301158 591658 301394
rect 591102 265158 591338 265394
rect 591422 265158 591658 265394
rect 591102 229158 591338 229394
rect 591422 229158 591658 229394
rect 591102 193158 591338 193394
rect 591422 193158 591658 193394
rect 591102 157158 591338 157394
rect 591422 157158 591658 157394
rect 591102 121158 591338 121394
rect 591422 121158 591658 121394
rect 591102 85158 591338 85394
rect 591422 85158 591658 85394
rect 591102 49158 591338 49394
rect 591422 49158 591658 49394
rect 591102 13158 591338 13394
rect 591422 13158 591658 13394
rect 591102 -6342 591338 -6106
rect 591422 -6342 591658 -6106
rect 591102 -6662 591338 -6426
rect 591422 -6662 591658 -6426
rect 592062 679158 592298 679394
rect 592382 679158 592618 679394
rect 592062 643158 592298 643394
rect 592382 643158 592618 643394
rect 592062 607158 592298 607394
rect 592382 607158 592618 607394
rect 592062 571158 592298 571394
rect 592382 571158 592618 571394
rect 592062 535158 592298 535394
rect 592382 535158 592618 535394
rect 592062 499158 592298 499394
rect 592382 499158 592618 499394
rect 592062 463158 592298 463394
rect 592382 463158 592618 463394
rect 592062 427158 592298 427394
rect 592382 427158 592618 427394
rect 592062 391158 592298 391394
rect 592382 391158 592618 391394
rect 592062 355158 592298 355394
rect 592382 355158 592618 355394
rect 592062 319158 592298 319394
rect 592382 319158 592618 319394
rect 592062 283158 592298 283394
rect 592382 283158 592618 283394
rect 592062 247158 592298 247394
rect 592382 247158 592618 247394
rect 592062 211158 592298 211394
rect 592382 211158 592618 211394
rect 592062 175158 592298 175394
rect 592382 175158 592618 175394
rect 592062 139158 592298 139394
rect 592382 139158 592618 139394
rect 592062 103158 592298 103394
rect 592382 103158 592618 103394
rect 592062 67158 592298 67394
rect 592382 67158 592618 67394
rect 592062 31158 592298 31394
rect 592382 31158 592618 31394
rect 570086 -7302 570322 -7066
rect 570086 -7622 570322 -7386
rect 592062 -7302 592298 -7066
rect 592382 -7302 592618 -7066
rect 592062 -7622 592298 -7386
rect 592382 -7622 592618 -7386
<< metal5 >>
rect -8726 711558 592650 711590
rect -8726 711322 -8694 711558
rect -8458 711322 -8374 711558
rect -8138 711322 30086 711558
rect 30322 711322 66086 711558
rect 66322 711322 102086 711558
rect 102322 711322 138086 711558
rect 138322 711322 174086 711558
rect 174322 711322 210086 711558
rect 210322 711322 246086 711558
rect 246322 711322 282086 711558
rect 282322 711322 318086 711558
rect 318322 711322 354086 711558
rect 354322 711322 390086 711558
rect 390322 711322 426086 711558
rect 426322 711322 462086 711558
rect 462322 711322 498086 711558
rect 498322 711322 534086 711558
rect 534322 711322 570086 711558
rect 570322 711322 592062 711558
rect 592298 711322 592382 711558
rect 592618 711322 592650 711558
rect -8726 711238 592650 711322
rect -8726 711002 -8694 711238
rect -8458 711002 -8374 711238
rect -8138 711002 30086 711238
rect 30322 711002 66086 711238
rect 66322 711002 102086 711238
rect 102322 711002 138086 711238
rect 138322 711002 174086 711238
rect 174322 711002 210086 711238
rect 210322 711002 246086 711238
rect 246322 711002 282086 711238
rect 282322 711002 318086 711238
rect 318322 711002 354086 711238
rect 354322 711002 390086 711238
rect 390322 711002 426086 711238
rect 426322 711002 462086 711238
rect 462322 711002 498086 711238
rect 498322 711002 534086 711238
rect 534322 711002 570086 711238
rect 570322 711002 592062 711238
rect 592298 711002 592382 711238
rect 592618 711002 592650 711238
rect -8726 710970 592650 711002
rect -7766 710598 591690 710630
rect -7766 710362 -7734 710598
rect -7498 710362 -7414 710598
rect -7178 710362 12086 710598
rect 12322 710362 48086 710598
rect 48322 710362 84086 710598
rect 84322 710362 120086 710598
rect 120322 710362 156086 710598
rect 156322 710362 192086 710598
rect 192322 710362 228086 710598
rect 228322 710362 264086 710598
rect 264322 710362 300086 710598
rect 300322 710362 336086 710598
rect 336322 710362 372086 710598
rect 372322 710362 408086 710598
rect 408322 710362 444086 710598
rect 444322 710362 480086 710598
rect 480322 710362 516086 710598
rect 516322 710362 552086 710598
rect 552322 710362 591102 710598
rect 591338 710362 591422 710598
rect 591658 710362 591690 710598
rect -7766 710278 591690 710362
rect -7766 710042 -7734 710278
rect -7498 710042 -7414 710278
rect -7178 710042 12086 710278
rect 12322 710042 48086 710278
rect 48322 710042 84086 710278
rect 84322 710042 120086 710278
rect 120322 710042 156086 710278
rect 156322 710042 192086 710278
rect 192322 710042 228086 710278
rect 228322 710042 264086 710278
rect 264322 710042 300086 710278
rect 300322 710042 336086 710278
rect 336322 710042 372086 710278
rect 372322 710042 408086 710278
rect 408322 710042 444086 710278
rect 444322 710042 480086 710278
rect 480322 710042 516086 710278
rect 516322 710042 552086 710278
rect 552322 710042 591102 710278
rect 591338 710042 591422 710278
rect 591658 710042 591690 710278
rect -7766 710010 591690 710042
rect -6806 709638 590730 709670
rect -6806 709402 -6774 709638
rect -6538 709402 -6454 709638
rect -6218 709402 26386 709638
rect 26622 709402 62386 709638
rect 62622 709402 98386 709638
rect 98622 709402 134386 709638
rect 134622 709402 170386 709638
rect 170622 709402 206386 709638
rect 206622 709402 242386 709638
rect 242622 709402 278386 709638
rect 278622 709402 314386 709638
rect 314622 709402 350386 709638
rect 350622 709402 386386 709638
rect 386622 709402 422386 709638
rect 422622 709402 458386 709638
rect 458622 709402 494386 709638
rect 494622 709402 530386 709638
rect 530622 709402 566386 709638
rect 566622 709402 590142 709638
rect 590378 709402 590462 709638
rect 590698 709402 590730 709638
rect -6806 709318 590730 709402
rect -6806 709082 -6774 709318
rect -6538 709082 -6454 709318
rect -6218 709082 26386 709318
rect 26622 709082 62386 709318
rect 62622 709082 98386 709318
rect 98622 709082 134386 709318
rect 134622 709082 170386 709318
rect 170622 709082 206386 709318
rect 206622 709082 242386 709318
rect 242622 709082 278386 709318
rect 278622 709082 314386 709318
rect 314622 709082 350386 709318
rect 350622 709082 386386 709318
rect 386622 709082 422386 709318
rect 422622 709082 458386 709318
rect 458622 709082 494386 709318
rect 494622 709082 530386 709318
rect 530622 709082 566386 709318
rect 566622 709082 590142 709318
rect 590378 709082 590462 709318
rect 590698 709082 590730 709318
rect -6806 709050 590730 709082
rect -5846 708678 589770 708710
rect -5846 708442 -5814 708678
rect -5578 708442 -5494 708678
rect -5258 708442 8386 708678
rect 8622 708442 44386 708678
rect 44622 708442 80386 708678
rect 80622 708442 116386 708678
rect 116622 708442 152386 708678
rect 152622 708442 188386 708678
rect 188622 708442 224386 708678
rect 224622 708442 260386 708678
rect 260622 708442 296386 708678
rect 296622 708442 332386 708678
rect 332622 708442 368386 708678
rect 368622 708442 404386 708678
rect 404622 708442 440386 708678
rect 440622 708442 476386 708678
rect 476622 708442 512386 708678
rect 512622 708442 548386 708678
rect 548622 708442 589182 708678
rect 589418 708442 589502 708678
rect 589738 708442 589770 708678
rect -5846 708358 589770 708442
rect -5846 708122 -5814 708358
rect -5578 708122 -5494 708358
rect -5258 708122 8386 708358
rect 8622 708122 44386 708358
rect 44622 708122 80386 708358
rect 80622 708122 116386 708358
rect 116622 708122 152386 708358
rect 152622 708122 188386 708358
rect 188622 708122 224386 708358
rect 224622 708122 260386 708358
rect 260622 708122 296386 708358
rect 296622 708122 332386 708358
rect 332622 708122 368386 708358
rect 368622 708122 404386 708358
rect 404622 708122 440386 708358
rect 440622 708122 476386 708358
rect 476622 708122 512386 708358
rect 512622 708122 548386 708358
rect 548622 708122 589182 708358
rect 589418 708122 589502 708358
rect 589738 708122 589770 708358
rect -5846 708090 589770 708122
rect -4886 707718 588810 707750
rect -4886 707482 -4854 707718
rect -4618 707482 -4534 707718
rect -4298 707482 22686 707718
rect 22922 707482 58686 707718
rect 58922 707482 94686 707718
rect 94922 707482 130686 707718
rect 130922 707482 166686 707718
rect 166922 707482 202686 707718
rect 202922 707482 238686 707718
rect 238922 707482 274686 707718
rect 274922 707482 310686 707718
rect 310922 707482 346686 707718
rect 346922 707482 382686 707718
rect 382922 707482 418686 707718
rect 418922 707482 454686 707718
rect 454922 707482 490686 707718
rect 490922 707482 526686 707718
rect 526922 707482 562686 707718
rect 562922 707482 588222 707718
rect 588458 707482 588542 707718
rect 588778 707482 588810 707718
rect -4886 707398 588810 707482
rect -4886 707162 -4854 707398
rect -4618 707162 -4534 707398
rect -4298 707162 22686 707398
rect 22922 707162 58686 707398
rect 58922 707162 94686 707398
rect 94922 707162 130686 707398
rect 130922 707162 166686 707398
rect 166922 707162 202686 707398
rect 202922 707162 238686 707398
rect 238922 707162 274686 707398
rect 274922 707162 310686 707398
rect 310922 707162 346686 707398
rect 346922 707162 382686 707398
rect 382922 707162 418686 707398
rect 418922 707162 454686 707398
rect 454922 707162 490686 707398
rect 490922 707162 526686 707398
rect 526922 707162 562686 707398
rect 562922 707162 588222 707398
rect 588458 707162 588542 707398
rect 588778 707162 588810 707398
rect -4886 707130 588810 707162
rect -3926 706758 587850 706790
rect -3926 706522 -3894 706758
rect -3658 706522 -3574 706758
rect -3338 706522 4686 706758
rect 4922 706522 40686 706758
rect 40922 706522 76686 706758
rect 76922 706522 112686 706758
rect 112922 706522 148686 706758
rect 148922 706522 184686 706758
rect 184922 706522 220686 706758
rect 220922 706522 256686 706758
rect 256922 706522 292686 706758
rect 292922 706522 328686 706758
rect 328922 706522 364686 706758
rect 364922 706522 400686 706758
rect 400922 706522 436686 706758
rect 436922 706522 472686 706758
rect 472922 706522 508686 706758
rect 508922 706522 544686 706758
rect 544922 706522 580686 706758
rect 580922 706522 587262 706758
rect 587498 706522 587582 706758
rect 587818 706522 587850 706758
rect -3926 706438 587850 706522
rect -3926 706202 -3894 706438
rect -3658 706202 -3574 706438
rect -3338 706202 4686 706438
rect 4922 706202 40686 706438
rect 40922 706202 76686 706438
rect 76922 706202 112686 706438
rect 112922 706202 148686 706438
rect 148922 706202 184686 706438
rect 184922 706202 220686 706438
rect 220922 706202 256686 706438
rect 256922 706202 292686 706438
rect 292922 706202 328686 706438
rect 328922 706202 364686 706438
rect 364922 706202 400686 706438
rect 400922 706202 436686 706438
rect 436922 706202 472686 706438
rect 472922 706202 508686 706438
rect 508922 706202 544686 706438
rect 544922 706202 580686 706438
rect 580922 706202 587262 706438
rect 587498 706202 587582 706438
rect 587818 706202 587850 706438
rect -3926 706170 587850 706202
rect -2966 705798 586890 705830
rect -2966 705562 -2934 705798
rect -2698 705562 -2614 705798
rect -2378 705562 18986 705798
rect 19222 705562 54986 705798
rect 55222 705562 90986 705798
rect 91222 705562 126986 705798
rect 127222 705562 162986 705798
rect 163222 705562 198986 705798
rect 199222 705562 234986 705798
rect 235222 705562 270986 705798
rect 271222 705562 306986 705798
rect 307222 705562 342986 705798
rect 343222 705562 378986 705798
rect 379222 705562 414986 705798
rect 415222 705562 450986 705798
rect 451222 705562 486986 705798
rect 487222 705562 522986 705798
rect 523222 705562 558986 705798
rect 559222 705562 586302 705798
rect 586538 705562 586622 705798
rect 586858 705562 586890 705798
rect -2966 705478 586890 705562
rect -2966 705242 -2934 705478
rect -2698 705242 -2614 705478
rect -2378 705242 18986 705478
rect 19222 705242 54986 705478
rect 55222 705242 90986 705478
rect 91222 705242 126986 705478
rect 127222 705242 162986 705478
rect 163222 705242 198986 705478
rect 199222 705242 234986 705478
rect 235222 705242 270986 705478
rect 271222 705242 306986 705478
rect 307222 705242 342986 705478
rect 343222 705242 378986 705478
rect 379222 705242 414986 705478
rect 415222 705242 450986 705478
rect 451222 705242 486986 705478
rect 487222 705242 522986 705478
rect 523222 705242 558986 705478
rect 559222 705242 586302 705478
rect 586538 705242 586622 705478
rect 586858 705242 586890 705478
rect -2966 705210 586890 705242
rect -2006 704838 585930 704870
rect -2006 704602 -1974 704838
rect -1738 704602 -1654 704838
rect -1418 704602 986 704838
rect 1222 704602 36986 704838
rect 37222 704602 72986 704838
rect 73222 704602 108986 704838
rect 109222 704602 144986 704838
rect 145222 704602 180986 704838
rect 181222 704602 216986 704838
rect 217222 704602 252986 704838
rect 253222 704602 288986 704838
rect 289222 704602 324986 704838
rect 325222 704602 360986 704838
rect 361222 704602 396986 704838
rect 397222 704602 432986 704838
rect 433222 704602 468986 704838
rect 469222 704602 504986 704838
rect 505222 704602 540986 704838
rect 541222 704602 576986 704838
rect 577222 704602 585342 704838
rect 585578 704602 585662 704838
rect 585898 704602 585930 704838
rect -2006 704518 585930 704602
rect -2006 704282 -1974 704518
rect -1738 704282 -1654 704518
rect -1418 704282 986 704518
rect 1222 704282 36986 704518
rect 37222 704282 72986 704518
rect 73222 704282 108986 704518
rect 109222 704282 144986 704518
rect 145222 704282 180986 704518
rect 181222 704282 216986 704518
rect 217222 704282 252986 704518
rect 253222 704282 288986 704518
rect 289222 704282 324986 704518
rect 325222 704282 360986 704518
rect 361222 704282 396986 704518
rect 397222 704282 432986 704518
rect 433222 704282 468986 704518
rect 469222 704282 504986 704518
rect 505222 704282 540986 704518
rect 541222 704282 576986 704518
rect 577222 704282 585342 704518
rect 585578 704282 585662 704518
rect 585898 704282 585930 704518
rect -2006 704250 585930 704282
rect -8726 697394 592650 697576
rect -8726 697158 -7734 697394
rect -7498 697158 -7414 697394
rect -7178 697158 12086 697394
rect 12322 697158 48086 697394
rect 48322 697158 84086 697394
rect 84322 697158 120086 697394
rect 120322 697158 156086 697394
rect 156322 697158 192086 697394
rect 192322 697158 228086 697394
rect 228322 697158 264086 697394
rect 264322 697158 300086 697394
rect 300322 697158 336086 697394
rect 336322 697158 372086 697394
rect 372322 697158 408086 697394
rect 408322 697158 444086 697394
rect 444322 697158 480086 697394
rect 480322 697158 516086 697394
rect 516322 697158 552086 697394
rect 552322 697158 591102 697394
rect 591338 697158 591422 697394
rect 591658 697158 592650 697394
rect -8726 696976 592650 697158
rect -6806 693694 590730 693876
rect -6806 693458 -5814 693694
rect -5578 693458 -5494 693694
rect -5258 693458 8386 693694
rect 8622 693458 44386 693694
rect 44622 693458 80386 693694
rect 80622 693458 116386 693694
rect 116622 693458 152386 693694
rect 152622 693458 188386 693694
rect 188622 693458 224386 693694
rect 224622 693458 260386 693694
rect 260622 693458 296386 693694
rect 296622 693458 332386 693694
rect 332622 693458 368386 693694
rect 368622 693458 404386 693694
rect 404622 693458 440386 693694
rect 440622 693458 476386 693694
rect 476622 693458 512386 693694
rect 512622 693458 548386 693694
rect 548622 693458 589182 693694
rect 589418 693458 589502 693694
rect 589738 693458 590730 693694
rect -6806 693276 590730 693458
rect -4886 689994 588810 690176
rect -4886 689758 -3894 689994
rect -3658 689758 -3574 689994
rect -3338 689758 4686 689994
rect 4922 689758 40686 689994
rect 40922 689758 76686 689994
rect 76922 689758 112686 689994
rect 112922 689758 148686 689994
rect 148922 689758 184686 689994
rect 184922 689758 220686 689994
rect 220922 689758 256686 689994
rect 256922 689758 292686 689994
rect 292922 689758 328686 689994
rect 328922 689758 364686 689994
rect 364922 689758 400686 689994
rect 400922 689758 436686 689994
rect 436922 689758 472686 689994
rect 472922 689758 508686 689994
rect 508922 689758 544686 689994
rect 544922 689758 580686 689994
rect 580922 689758 587262 689994
rect 587498 689758 587582 689994
rect 587818 689758 588810 689994
rect -4886 689576 588810 689758
rect -2966 686294 586890 686476
rect -2966 686058 -1974 686294
rect -1738 686058 -1654 686294
rect -1418 686058 986 686294
rect 1222 686058 36986 686294
rect 37222 686058 72986 686294
rect 73222 686058 108986 686294
rect 109222 686058 144986 686294
rect 145222 686058 180986 686294
rect 181222 686058 216986 686294
rect 217222 686058 252986 686294
rect 253222 686058 288986 686294
rect 289222 686058 324986 686294
rect 325222 686058 360986 686294
rect 361222 686058 396986 686294
rect 397222 686058 432986 686294
rect 433222 686058 468986 686294
rect 469222 686058 504986 686294
rect 505222 686058 540986 686294
rect 541222 686058 576986 686294
rect 577222 686058 585342 686294
rect 585578 686058 585662 686294
rect 585898 686058 586890 686294
rect -2966 685876 586890 686058
rect -8726 679394 592650 679576
rect -8726 679158 -8694 679394
rect -8458 679158 -8374 679394
rect -8138 679158 30086 679394
rect 30322 679158 66086 679394
rect 66322 679158 102086 679394
rect 102322 679158 138086 679394
rect 138322 679158 174086 679394
rect 174322 679158 210086 679394
rect 210322 679158 246086 679394
rect 246322 679158 282086 679394
rect 282322 679158 318086 679394
rect 318322 679158 354086 679394
rect 354322 679158 390086 679394
rect 390322 679158 426086 679394
rect 426322 679158 462086 679394
rect 462322 679158 498086 679394
rect 498322 679158 534086 679394
rect 534322 679158 570086 679394
rect 570322 679158 592062 679394
rect 592298 679158 592382 679394
rect 592618 679158 592650 679394
rect -8726 678976 592650 679158
rect -6806 675694 590730 675876
rect -6806 675458 -6774 675694
rect -6538 675458 -6454 675694
rect -6218 675458 26386 675694
rect 26622 675458 62386 675694
rect 62622 675458 98386 675694
rect 98622 675458 134386 675694
rect 134622 675458 170386 675694
rect 170622 675458 206386 675694
rect 206622 675458 242386 675694
rect 242622 675458 278386 675694
rect 278622 675458 314386 675694
rect 314622 675458 350386 675694
rect 350622 675458 386386 675694
rect 386622 675458 422386 675694
rect 422622 675458 458386 675694
rect 458622 675458 494386 675694
rect 494622 675458 530386 675694
rect 530622 675458 566386 675694
rect 566622 675458 590142 675694
rect 590378 675458 590462 675694
rect 590698 675458 590730 675694
rect -6806 675276 590730 675458
rect -4886 671994 588810 672176
rect -4886 671758 -4854 671994
rect -4618 671758 -4534 671994
rect -4298 671758 22686 671994
rect 22922 671758 58686 671994
rect 58922 671758 94686 671994
rect 94922 671758 130686 671994
rect 130922 671758 166686 671994
rect 166922 671758 202686 671994
rect 202922 671758 238686 671994
rect 238922 671758 274686 671994
rect 274922 671758 310686 671994
rect 310922 671758 346686 671994
rect 346922 671758 382686 671994
rect 382922 671758 418686 671994
rect 418922 671758 454686 671994
rect 454922 671758 490686 671994
rect 490922 671758 526686 671994
rect 526922 671758 562686 671994
rect 562922 671758 588222 671994
rect 588458 671758 588542 671994
rect 588778 671758 588810 671994
rect -4886 671576 588810 671758
rect -2966 668294 586890 668476
rect -2966 668058 -2934 668294
rect -2698 668058 -2614 668294
rect -2378 668058 18986 668294
rect 19222 668058 54986 668294
rect 55222 668058 90986 668294
rect 91222 668058 126986 668294
rect 127222 668058 162986 668294
rect 163222 668058 198986 668294
rect 199222 668058 234986 668294
rect 235222 668058 270986 668294
rect 271222 668058 306986 668294
rect 307222 668058 342986 668294
rect 343222 668058 378986 668294
rect 379222 668058 414986 668294
rect 415222 668058 450986 668294
rect 451222 668058 486986 668294
rect 487222 668058 522986 668294
rect 523222 668058 558986 668294
rect 559222 668058 586302 668294
rect 586538 668058 586622 668294
rect 586858 668058 586890 668294
rect -2966 667876 586890 668058
rect -8726 661394 592650 661576
rect -8726 661158 -7734 661394
rect -7498 661158 -7414 661394
rect -7178 661158 12086 661394
rect 12322 661158 48086 661394
rect 48322 661158 84086 661394
rect 84322 661158 120086 661394
rect 120322 661158 156086 661394
rect 156322 661158 192086 661394
rect 192322 661158 228086 661394
rect 228322 661158 264086 661394
rect 264322 661158 300086 661394
rect 300322 661158 336086 661394
rect 336322 661158 372086 661394
rect 372322 661158 408086 661394
rect 408322 661158 444086 661394
rect 444322 661158 480086 661394
rect 480322 661158 516086 661394
rect 516322 661158 552086 661394
rect 552322 661158 591102 661394
rect 591338 661158 591422 661394
rect 591658 661158 592650 661394
rect -8726 660976 592650 661158
rect -6806 657694 590730 657876
rect -6806 657458 -5814 657694
rect -5578 657458 -5494 657694
rect -5258 657458 8386 657694
rect 8622 657458 44386 657694
rect 44622 657458 80386 657694
rect 80622 657458 116386 657694
rect 116622 657458 152386 657694
rect 152622 657458 188386 657694
rect 188622 657458 224386 657694
rect 224622 657458 260386 657694
rect 260622 657458 296386 657694
rect 296622 657458 332386 657694
rect 332622 657458 368386 657694
rect 368622 657458 404386 657694
rect 404622 657458 440386 657694
rect 440622 657458 476386 657694
rect 476622 657458 512386 657694
rect 512622 657458 548386 657694
rect 548622 657458 589182 657694
rect 589418 657458 589502 657694
rect 589738 657458 590730 657694
rect -6806 657276 590730 657458
rect -4886 653994 588810 654176
rect -4886 653758 -3894 653994
rect -3658 653758 -3574 653994
rect -3338 653758 4686 653994
rect 4922 653758 40686 653994
rect 40922 653758 76686 653994
rect 76922 653758 112686 653994
rect 112922 653758 148686 653994
rect 148922 653758 184686 653994
rect 184922 653758 220686 653994
rect 220922 653758 256686 653994
rect 256922 653758 292686 653994
rect 292922 653758 328686 653994
rect 328922 653758 364686 653994
rect 364922 653758 400686 653994
rect 400922 653758 436686 653994
rect 436922 653758 472686 653994
rect 472922 653758 508686 653994
rect 508922 653758 544686 653994
rect 544922 653758 580686 653994
rect 580922 653758 587262 653994
rect 587498 653758 587582 653994
rect 587818 653758 588810 653994
rect -4886 653576 588810 653758
rect -2966 650294 586890 650476
rect -2966 650058 -1974 650294
rect -1738 650058 -1654 650294
rect -1418 650058 986 650294
rect 1222 650058 36986 650294
rect 37222 650058 72986 650294
rect 73222 650058 108986 650294
rect 109222 650058 144986 650294
rect 145222 650058 180986 650294
rect 181222 650058 216986 650294
rect 217222 650058 252986 650294
rect 253222 650058 288986 650294
rect 289222 650058 324986 650294
rect 325222 650058 360986 650294
rect 361222 650058 396986 650294
rect 397222 650058 432986 650294
rect 433222 650058 468986 650294
rect 469222 650058 504986 650294
rect 505222 650058 540986 650294
rect 541222 650058 576986 650294
rect 577222 650058 585342 650294
rect 585578 650058 585662 650294
rect 585898 650058 586890 650294
rect -2966 649876 586890 650058
rect -8726 643394 592650 643576
rect -8726 643158 -8694 643394
rect -8458 643158 -8374 643394
rect -8138 643158 30086 643394
rect 30322 643158 66086 643394
rect 66322 643158 102086 643394
rect 102322 643158 138086 643394
rect 138322 643158 174086 643394
rect 174322 643158 210086 643394
rect 210322 643158 246086 643394
rect 246322 643158 282086 643394
rect 282322 643158 318086 643394
rect 318322 643158 354086 643394
rect 354322 643158 390086 643394
rect 390322 643158 426086 643394
rect 426322 643158 462086 643394
rect 462322 643158 498086 643394
rect 498322 643158 534086 643394
rect 534322 643158 570086 643394
rect 570322 643158 592062 643394
rect 592298 643158 592382 643394
rect 592618 643158 592650 643394
rect -8726 642976 592650 643158
rect -6806 639694 590730 639876
rect -6806 639458 -6774 639694
rect -6538 639458 -6454 639694
rect -6218 639458 26386 639694
rect 26622 639458 62386 639694
rect 62622 639458 98386 639694
rect 98622 639458 134386 639694
rect 134622 639458 170386 639694
rect 170622 639458 206386 639694
rect 206622 639458 242386 639694
rect 242622 639458 278386 639694
rect 278622 639458 314386 639694
rect 314622 639458 350386 639694
rect 350622 639458 386386 639694
rect 386622 639458 422386 639694
rect 422622 639458 458386 639694
rect 458622 639458 494386 639694
rect 494622 639458 530386 639694
rect 530622 639458 566386 639694
rect 566622 639458 590142 639694
rect 590378 639458 590462 639694
rect 590698 639458 590730 639694
rect -6806 639276 590730 639458
rect -4886 635994 588810 636176
rect -4886 635758 -4854 635994
rect -4618 635758 -4534 635994
rect -4298 635758 22686 635994
rect 22922 635758 58686 635994
rect 58922 635758 94686 635994
rect 94922 635758 130686 635994
rect 130922 635758 166686 635994
rect 166922 635758 202686 635994
rect 202922 635758 238686 635994
rect 238922 635758 274686 635994
rect 274922 635758 310686 635994
rect 310922 635758 346686 635994
rect 346922 635758 382686 635994
rect 382922 635758 418686 635994
rect 418922 635758 454686 635994
rect 454922 635758 490686 635994
rect 490922 635758 526686 635994
rect 526922 635758 562686 635994
rect 562922 635758 588222 635994
rect 588458 635758 588542 635994
rect 588778 635758 588810 635994
rect -4886 635576 588810 635758
rect -2966 632294 586890 632476
rect -2966 632058 -2934 632294
rect -2698 632058 -2614 632294
rect -2378 632058 18986 632294
rect 19222 632058 54986 632294
rect 55222 632058 90986 632294
rect 91222 632058 126986 632294
rect 127222 632058 162986 632294
rect 163222 632058 198986 632294
rect 199222 632058 234986 632294
rect 235222 632058 270986 632294
rect 271222 632058 306986 632294
rect 307222 632058 342986 632294
rect 343222 632058 378986 632294
rect 379222 632058 414986 632294
rect 415222 632058 450986 632294
rect 451222 632058 486986 632294
rect 487222 632058 522986 632294
rect 523222 632058 558986 632294
rect 559222 632058 586302 632294
rect 586538 632058 586622 632294
rect 586858 632058 586890 632294
rect -2966 631876 586890 632058
rect -8726 625394 592650 625576
rect -8726 625158 -7734 625394
rect -7498 625158 -7414 625394
rect -7178 625158 12086 625394
rect 12322 625158 48086 625394
rect 48322 625158 84086 625394
rect 84322 625158 120086 625394
rect 120322 625158 156086 625394
rect 156322 625158 192086 625394
rect 192322 625158 228086 625394
rect 228322 625158 264086 625394
rect 264322 625158 300086 625394
rect 300322 625158 336086 625394
rect 336322 625158 372086 625394
rect 372322 625158 408086 625394
rect 408322 625158 444086 625394
rect 444322 625158 480086 625394
rect 480322 625158 516086 625394
rect 516322 625158 552086 625394
rect 552322 625158 591102 625394
rect 591338 625158 591422 625394
rect 591658 625158 592650 625394
rect -8726 624976 592650 625158
rect -6806 621694 590730 621876
rect -6806 621458 -5814 621694
rect -5578 621458 -5494 621694
rect -5258 621458 8386 621694
rect 8622 621458 44386 621694
rect 44622 621458 80386 621694
rect 80622 621458 116386 621694
rect 116622 621458 152386 621694
rect 152622 621458 188386 621694
rect 188622 621458 224386 621694
rect 224622 621458 260386 621694
rect 260622 621458 296386 621694
rect 296622 621458 332386 621694
rect 332622 621458 368386 621694
rect 368622 621458 404386 621694
rect 404622 621458 440386 621694
rect 440622 621458 476386 621694
rect 476622 621458 512386 621694
rect 512622 621458 548386 621694
rect 548622 621458 589182 621694
rect 589418 621458 589502 621694
rect 589738 621458 590730 621694
rect -6806 621276 590730 621458
rect -4886 617994 588810 618176
rect -4886 617758 -3894 617994
rect -3658 617758 -3574 617994
rect -3338 617758 4686 617994
rect 4922 617758 40686 617994
rect 40922 617758 76686 617994
rect 76922 617758 112686 617994
rect 112922 617758 148686 617994
rect 148922 617758 184686 617994
rect 184922 617758 220686 617994
rect 220922 617758 256686 617994
rect 256922 617758 292686 617994
rect 292922 617758 328686 617994
rect 328922 617758 364686 617994
rect 364922 617758 400686 617994
rect 400922 617758 436686 617994
rect 436922 617758 472686 617994
rect 472922 617758 508686 617994
rect 508922 617758 544686 617994
rect 544922 617758 580686 617994
rect 580922 617758 587262 617994
rect 587498 617758 587582 617994
rect 587818 617758 588810 617994
rect -4886 617576 588810 617758
rect -2966 614294 586890 614476
rect -2966 614058 -1974 614294
rect -1738 614058 -1654 614294
rect -1418 614058 986 614294
rect 1222 614058 36986 614294
rect 37222 614058 72986 614294
rect 73222 614058 108986 614294
rect 109222 614058 144986 614294
rect 145222 614058 180986 614294
rect 181222 614058 216986 614294
rect 217222 614058 252986 614294
rect 253222 614058 288986 614294
rect 289222 614058 324986 614294
rect 325222 614058 360986 614294
rect 361222 614058 396986 614294
rect 397222 614058 432986 614294
rect 433222 614058 468986 614294
rect 469222 614058 504986 614294
rect 505222 614058 540986 614294
rect 541222 614058 576986 614294
rect 577222 614058 585342 614294
rect 585578 614058 585662 614294
rect 585898 614058 586890 614294
rect -2966 613876 586890 614058
rect -8726 607394 592650 607576
rect -8726 607158 -8694 607394
rect -8458 607158 -8374 607394
rect -8138 607158 30086 607394
rect 30322 607158 66086 607394
rect 66322 607158 102086 607394
rect 102322 607158 138086 607394
rect 138322 607158 174086 607394
rect 174322 607158 210086 607394
rect 210322 607158 246086 607394
rect 246322 607158 282086 607394
rect 282322 607158 318086 607394
rect 318322 607158 354086 607394
rect 354322 607158 390086 607394
rect 390322 607158 426086 607394
rect 426322 607158 462086 607394
rect 462322 607158 498086 607394
rect 498322 607158 534086 607394
rect 534322 607158 570086 607394
rect 570322 607158 592062 607394
rect 592298 607158 592382 607394
rect 592618 607158 592650 607394
rect -8726 606976 592650 607158
rect -6806 603694 590730 603876
rect -6806 603458 -6774 603694
rect -6538 603458 -6454 603694
rect -6218 603458 26386 603694
rect 26622 603458 62386 603694
rect 62622 603458 98386 603694
rect 98622 603458 134386 603694
rect 134622 603458 170386 603694
rect 170622 603458 206386 603694
rect 206622 603458 242386 603694
rect 242622 603458 278386 603694
rect 278622 603458 314386 603694
rect 314622 603458 350386 603694
rect 350622 603458 386386 603694
rect 386622 603458 422386 603694
rect 422622 603458 458386 603694
rect 458622 603458 494386 603694
rect 494622 603458 530386 603694
rect 530622 603458 566386 603694
rect 566622 603458 590142 603694
rect 590378 603458 590462 603694
rect 590698 603458 590730 603694
rect -6806 603276 590730 603458
rect -4886 599994 588810 600176
rect -4886 599758 -4854 599994
rect -4618 599758 -4534 599994
rect -4298 599758 22686 599994
rect 22922 599758 58686 599994
rect 58922 599758 94686 599994
rect 94922 599758 130686 599994
rect 130922 599758 166686 599994
rect 166922 599758 202686 599994
rect 202922 599758 238686 599994
rect 238922 599758 274686 599994
rect 274922 599758 310686 599994
rect 310922 599758 346686 599994
rect 346922 599758 382686 599994
rect 382922 599758 418686 599994
rect 418922 599758 454686 599994
rect 454922 599758 490686 599994
rect 490922 599758 526686 599994
rect 526922 599758 562686 599994
rect 562922 599758 588222 599994
rect 588458 599758 588542 599994
rect 588778 599758 588810 599994
rect -4886 599576 588810 599758
rect -2966 596294 586890 596476
rect -2966 596058 -2934 596294
rect -2698 596058 -2614 596294
rect -2378 596058 18986 596294
rect 19222 596058 54986 596294
rect 55222 596058 90986 596294
rect 91222 596058 126986 596294
rect 127222 596058 162986 596294
rect 163222 596058 198986 596294
rect 199222 596058 234986 596294
rect 235222 596058 270986 596294
rect 271222 596058 306986 596294
rect 307222 596058 342986 596294
rect 343222 596058 378986 596294
rect 379222 596058 414986 596294
rect 415222 596058 450986 596294
rect 451222 596058 486986 596294
rect 487222 596058 522986 596294
rect 523222 596058 558986 596294
rect 559222 596058 586302 596294
rect 586538 596058 586622 596294
rect 586858 596058 586890 596294
rect -2966 595876 586890 596058
rect -8726 589394 592650 589576
rect -8726 589158 -7734 589394
rect -7498 589158 -7414 589394
rect -7178 589158 12086 589394
rect 12322 589158 48086 589394
rect 48322 589158 84086 589394
rect 84322 589158 120086 589394
rect 120322 589158 156086 589394
rect 156322 589158 192086 589394
rect 192322 589158 228086 589394
rect 228322 589158 264086 589394
rect 264322 589158 300086 589394
rect 300322 589158 336086 589394
rect 336322 589158 372086 589394
rect 372322 589158 408086 589394
rect 408322 589158 444086 589394
rect 444322 589158 480086 589394
rect 480322 589158 516086 589394
rect 516322 589158 552086 589394
rect 552322 589158 591102 589394
rect 591338 589158 591422 589394
rect 591658 589158 592650 589394
rect -8726 588976 592650 589158
rect -6806 585694 590730 585876
rect -6806 585458 -5814 585694
rect -5578 585458 -5494 585694
rect -5258 585458 8386 585694
rect 8622 585458 44386 585694
rect 44622 585458 80386 585694
rect 80622 585458 116386 585694
rect 116622 585458 152386 585694
rect 152622 585458 188386 585694
rect 188622 585458 224386 585694
rect 224622 585458 260386 585694
rect 260622 585458 296386 585694
rect 296622 585458 332386 585694
rect 332622 585458 368386 585694
rect 368622 585458 404386 585694
rect 404622 585458 440386 585694
rect 440622 585458 476386 585694
rect 476622 585458 512386 585694
rect 512622 585458 548386 585694
rect 548622 585458 589182 585694
rect 589418 585458 589502 585694
rect 589738 585458 590730 585694
rect -6806 585276 590730 585458
rect -4886 581994 588810 582176
rect -4886 581758 -3894 581994
rect -3658 581758 -3574 581994
rect -3338 581758 4686 581994
rect 4922 581758 40686 581994
rect 40922 581758 76686 581994
rect 76922 581758 112686 581994
rect 112922 581758 148686 581994
rect 148922 581758 184686 581994
rect 184922 581758 220686 581994
rect 220922 581758 256686 581994
rect 256922 581758 292686 581994
rect 292922 581758 328686 581994
rect 328922 581758 364686 581994
rect 364922 581758 400686 581994
rect 400922 581758 436686 581994
rect 436922 581758 472686 581994
rect 472922 581758 508686 581994
rect 508922 581758 544686 581994
rect 544922 581758 580686 581994
rect 580922 581758 587262 581994
rect 587498 581758 587582 581994
rect 587818 581758 588810 581994
rect -4886 581576 588810 581758
rect -2966 578294 586890 578476
rect -2966 578058 -1974 578294
rect -1738 578058 -1654 578294
rect -1418 578058 986 578294
rect 1222 578058 36986 578294
rect 37222 578058 72986 578294
rect 73222 578058 108986 578294
rect 109222 578058 144986 578294
rect 145222 578058 180986 578294
rect 181222 578058 216986 578294
rect 217222 578058 252986 578294
rect 253222 578058 288986 578294
rect 289222 578058 324986 578294
rect 325222 578058 360986 578294
rect 361222 578058 396986 578294
rect 397222 578058 432986 578294
rect 433222 578058 468986 578294
rect 469222 578058 504986 578294
rect 505222 578058 540986 578294
rect 541222 578058 576986 578294
rect 577222 578058 585342 578294
rect 585578 578058 585662 578294
rect 585898 578058 586890 578294
rect -2966 577876 586890 578058
rect -8726 571394 592650 571576
rect -8726 571158 -8694 571394
rect -8458 571158 -8374 571394
rect -8138 571158 30086 571394
rect 30322 571158 66086 571394
rect 66322 571158 102086 571394
rect 102322 571158 138086 571394
rect 138322 571158 174086 571394
rect 174322 571158 210086 571394
rect 210322 571158 246086 571394
rect 246322 571158 282086 571394
rect 282322 571158 318086 571394
rect 318322 571158 354086 571394
rect 354322 571158 390086 571394
rect 390322 571158 426086 571394
rect 426322 571158 462086 571394
rect 462322 571158 498086 571394
rect 498322 571158 534086 571394
rect 534322 571158 570086 571394
rect 570322 571158 592062 571394
rect 592298 571158 592382 571394
rect 592618 571158 592650 571394
rect -8726 570976 592650 571158
rect -6806 567694 590730 567876
rect -6806 567458 -6774 567694
rect -6538 567458 -6454 567694
rect -6218 567458 26386 567694
rect 26622 567458 62386 567694
rect 62622 567458 98386 567694
rect 98622 567458 134386 567694
rect 134622 567458 170386 567694
rect 170622 567458 206386 567694
rect 206622 567458 242386 567694
rect 242622 567458 278386 567694
rect 278622 567458 314386 567694
rect 314622 567458 350386 567694
rect 350622 567458 386386 567694
rect 386622 567458 422386 567694
rect 422622 567458 458386 567694
rect 458622 567458 494386 567694
rect 494622 567458 530386 567694
rect 530622 567458 566386 567694
rect 566622 567458 590142 567694
rect 590378 567458 590462 567694
rect 590698 567458 590730 567694
rect -6806 567276 590730 567458
rect -4886 563994 588810 564176
rect -4886 563758 -4854 563994
rect -4618 563758 -4534 563994
rect -4298 563758 22686 563994
rect 22922 563758 58686 563994
rect 58922 563758 94686 563994
rect 94922 563758 130686 563994
rect 130922 563758 166686 563994
rect 166922 563758 202686 563994
rect 202922 563758 238686 563994
rect 238922 563758 274686 563994
rect 274922 563758 310686 563994
rect 310922 563758 346686 563994
rect 346922 563758 382686 563994
rect 382922 563758 418686 563994
rect 418922 563758 454686 563994
rect 454922 563758 490686 563994
rect 490922 563758 526686 563994
rect 526922 563758 562686 563994
rect 562922 563758 588222 563994
rect 588458 563758 588542 563994
rect 588778 563758 588810 563994
rect -4886 563576 588810 563758
rect -2966 560294 586890 560476
rect -2966 560058 -2934 560294
rect -2698 560058 -2614 560294
rect -2378 560058 18986 560294
rect 19222 560058 54986 560294
rect 55222 560058 90986 560294
rect 91222 560058 126986 560294
rect 127222 560058 162986 560294
rect 163222 560058 198986 560294
rect 199222 560058 234986 560294
rect 235222 560058 270986 560294
rect 271222 560058 306986 560294
rect 307222 560058 342986 560294
rect 343222 560058 378986 560294
rect 379222 560058 414986 560294
rect 415222 560058 450986 560294
rect 451222 560058 486986 560294
rect 487222 560058 522986 560294
rect 523222 560058 558986 560294
rect 559222 560058 586302 560294
rect 586538 560058 586622 560294
rect 586858 560058 586890 560294
rect -2966 559876 586890 560058
rect -8726 553394 592650 553576
rect -8726 553158 -7734 553394
rect -7498 553158 -7414 553394
rect -7178 553158 12086 553394
rect 12322 553158 48086 553394
rect 48322 553158 84086 553394
rect 84322 553158 120086 553394
rect 120322 553158 156086 553394
rect 156322 553158 192086 553394
rect 192322 553158 228086 553394
rect 228322 553158 264086 553394
rect 264322 553158 300086 553394
rect 300322 553158 336086 553394
rect 336322 553158 372086 553394
rect 372322 553158 408086 553394
rect 408322 553158 444086 553394
rect 444322 553158 480086 553394
rect 480322 553158 516086 553394
rect 516322 553158 552086 553394
rect 552322 553158 591102 553394
rect 591338 553158 591422 553394
rect 591658 553158 592650 553394
rect -8726 552976 592650 553158
rect -6806 549694 590730 549876
rect -6806 549458 -5814 549694
rect -5578 549458 -5494 549694
rect -5258 549458 8386 549694
rect 8622 549458 44386 549694
rect 44622 549458 80386 549694
rect 80622 549458 116386 549694
rect 116622 549458 152386 549694
rect 152622 549458 188386 549694
rect 188622 549458 224386 549694
rect 224622 549458 260386 549694
rect 260622 549458 296386 549694
rect 296622 549458 332386 549694
rect 332622 549458 368386 549694
rect 368622 549458 404386 549694
rect 404622 549458 440386 549694
rect 440622 549458 476386 549694
rect 476622 549458 512386 549694
rect 512622 549458 548386 549694
rect 548622 549458 589182 549694
rect 589418 549458 589502 549694
rect 589738 549458 590730 549694
rect -6806 549276 590730 549458
rect -4886 545994 588810 546176
rect -4886 545758 -3894 545994
rect -3658 545758 -3574 545994
rect -3338 545758 4686 545994
rect 4922 545758 40686 545994
rect 40922 545758 76686 545994
rect 76922 545758 112686 545994
rect 112922 545758 148686 545994
rect 148922 545758 184686 545994
rect 184922 545758 220686 545994
rect 220922 545758 256686 545994
rect 256922 545758 292686 545994
rect 292922 545758 328686 545994
rect 328922 545758 364686 545994
rect 364922 545758 400686 545994
rect 400922 545758 436686 545994
rect 436922 545758 472686 545994
rect 472922 545758 508686 545994
rect 508922 545758 544686 545994
rect 544922 545758 580686 545994
rect 580922 545758 587262 545994
rect 587498 545758 587582 545994
rect 587818 545758 588810 545994
rect -4886 545576 588810 545758
rect -2966 542294 586890 542476
rect -2966 542058 -1974 542294
rect -1738 542058 -1654 542294
rect -1418 542058 986 542294
rect 1222 542058 36986 542294
rect 37222 542058 72986 542294
rect 73222 542058 108986 542294
rect 109222 542058 144986 542294
rect 145222 542058 180986 542294
rect 181222 542058 216986 542294
rect 217222 542058 252986 542294
rect 253222 542058 288986 542294
rect 289222 542058 324986 542294
rect 325222 542058 360986 542294
rect 361222 542058 396986 542294
rect 397222 542058 432986 542294
rect 433222 542058 468986 542294
rect 469222 542058 504986 542294
rect 505222 542058 540986 542294
rect 541222 542058 576986 542294
rect 577222 542058 585342 542294
rect 585578 542058 585662 542294
rect 585898 542058 586890 542294
rect -2966 541876 586890 542058
rect -8726 535394 592650 535576
rect -8726 535158 -8694 535394
rect -8458 535158 -8374 535394
rect -8138 535158 30086 535394
rect 30322 535158 66086 535394
rect 66322 535158 102086 535394
rect 102322 535158 138086 535394
rect 138322 535158 174086 535394
rect 174322 535158 210086 535394
rect 210322 535158 246086 535394
rect 246322 535158 282086 535394
rect 282322 535158 318086 535394
rect 318322 535158 354086 535394
rect 354322 535158 390086 535394
rect 390322 535158 426086 535394
rect 426322 535158 462086 535394
rect 462322 535158 498086 535394
rect 498322 535158 534086 535394
rect 534322 535158 570086 535394
rect 570322 535158 592062 535394
rect 592298 535158 592382 535394
rect 592618 535158 592650 535394
rect -8726 534976 592650 535158
rect -6806 531694 590730 531876
rect -6806 531458 -6774 531694
rect -6538 531458 -6454 531694
rect -6218 531458 26386 531694
rect 26622 531458 62386 531694
rect 62622 531458 98386 531694
rect 98622 531458 134386 531694
rect 134622 531458 170386 531694
rect 170622 531458 206386 531694
rect 206622 531458 242386 531694
rect 242622 531458 278386 531694
rect 278622 531458 314386 531694
rect 314622 531458 350386 531694
rect 350622 531458 386386 531694
rect 386622 531458 422386 531694
rect 422622 531458 458386 531694
rect 458622 531458 494386 531694
rect 494622 531458 530386 531694
rect 530622 531458 566386 531694
rect 566622 531458 590142 531694
rect 590378 531458 590462 531694
rect 590698 531458 590730 531694
rect -6806 531276 590730 531458
rect -4886 527994 588810 528176
rect -4886 527758 -4854 527994
rect -4618 527758 -4534 527994
rect -4298 527758 22686 527994
rect 22922 527758 58686 527994
rect 58922 527758 94686 527994
rect 94922 527758 130686 527994
rect 130922 527758 166686 527994
rect 166922 527758 202686 527994
rect 202922 527758 238686 527994
rect 238922 527758 274686 527994
rect 274922 527758 310686 527994
rect 310922 527758 346686 527994
rect 346922 527758 382686 527994
rect 382922 527758 418686 527994
rect 418922 527758 454686 527994
rect 454922 527758 490686 527994
rect 490922 527758 526686 527994
rect 526922 527758 562686 527994
rect 562922 527758 588222 527994
rect 588458 527758 588542 527994
rect 588778 527758 588810 527994
rect -4886 527576 588810 527758
rect -2966 524294 586890 524476
rect -2966 524058 -2934 524294
rect -2698 524058 -2614 524294
rect -2378 524058 18986 524294
rect 19222 524058 54986 524294
rect 55222 524058 90986 524294
rect 91222 524058 126986 524294
rect 127222 524058 162986 524294
rect 163222 524058 198986 524294
rect 199222 524058 234986 524294
rect 235222 524058 270986 524294
rect 271222 524058 306986 524294
rect 307222 524058 342986 524294
rect 343222 524058 378986 524294
rect 379222 524058 414986 524294
rect 415222 524058 450986 524294
rect 451222 524058 486986 524294
rect 487222 524058 522986 524294
rect 523222 524058 558986 524294
rect 559222 524058 586302 524294
rect 586538 524058 586622 524294
rect 586858 524058 586890 524294
rect -2966 523876 586890 524058
rect -8726 517394 592650 517576
rect -8726 517158 -7734 517394
rect -7498 517158 -7414 517394
rect -7178 517158 12086 517394
rect 12322 517158 48086 517394
rect 48322 517158 84086 517394
rect 84322 517158 120086 517394
rect 120322 517158 156086 517394
rect 156322 517158 192086 517394
rect 192322 517158 228086 517394
rect 228322 517158 264086 517394
rect 264322 517158 300086 517394
rect 300322 517158 336086 517394
rect 336322 517158 372086 517394
rect 372322 517158 408086 517394
rect 408322 517158 444086 517394
rect 444322 517158 480086 517394
rect 480322 517158 516086 517394
rect 516322 517158 552086 517394
rect 552322 517158 591102 517394
rect 591338 517158 591422 517394
rect 591658 517158 592650 517394
rect -8726 516976 592650 517158
rect -6806 513694 590730 513876
rect -6806 513458 -5814 513694
rect -5578 513458 -5494 513694
rect -5258 513458 8386 513694
rect 8622 513458 44386 513694
rect 44622 513458 80386 513694
rect 80622 513458 116386 513694
rect 116622 513458 152386 513694
rect 152622 513458 188386 513694
rect 188622 513458 224386 513694
rect 224622 513458 260386 513694
rect 260622 513458 296386 513694
rect 296622 513458 332386 513694
rect 332622 513458 368386 513694
rect 368622 513458 404386 513694
rect 404622 513458 440386 513694
rect 440622 513458 476386 513694
rect 476622 513458 512386 513694
rect 512622 513458 548386 513694
rect 548622 513458 589182 513694
rect 589418 513458 589502 513694
rect 589738 513458 590730 513694
rect -6806 513276 590730 513458
rect -4886 509994 588810 510176
rect -4886 509758 -3894 509994
rect -3658 509758 -3574 509994
rect -3338 509758 4686 509994
rect 4922 509758 40686 509994
rect 40922 509758 76686 509994
rect 76922 509758 112686 509994
rect 112922 509758 148686 509994
rect 148922 509758 184686 509994
rect 184922 509758 220686 509994
rect 220922 509758 256686 509994
rect 256922 509758 292686 509994
rect 292922 509758 328686 509994
rect 328922 509758 364686 509994
rect 364922 509758 400686 509994
rect 400922 509758 436686 509994
rect 436922 509758 472686 509994
rect 472922 509758 508686 509994
rect 508922 509758 544686 509994
rect 544922 509758 580686 509994
rect 580922 509758 587262 509994
rect 587498 509758 587582 509994
rect 587818 509758 588810 509994
rect -4886 509576 588810 509758
rect -2966 506294 586890 506476
rect -2966 506058 -1974 506294
rect -1738 506058 -1654 506294
rect -1418 506058 986 506294
rect 1222 506058 36986 506294
rect 37222 506058 72986 506294
rect 73222 506058 108986 506294
rect 109222 506058 144986 506294
rect 145222 506058 180986 506294
rect 181222 506058 216986 506294
rect 217222 506058 252986 506294
rect 253222 506058 288986 506294
rect 289222 506058 324986 506294
rect 325222 506058 360986 506294
rect 361222 506058 396986 506294
rect 397222 506058 432986 506294
rect 433222 506058 468986 506294
rect 469222 506058 504986 506294
rect 505222 506058 540986 506294
rect 541222 506058 576986 506294
rect 577222 506058 585342 506294
rect 585578 506058 585662 506294
rect 585898 506058 586890 506294
rect -2966 505876 586890 506058
rect -8726 499394 592650 499576
rect -8726 499158 -8694 499394
rect -8458 499158 -8374 499394
rect -8138 499158 30086 499394
rect 30322 499158 66086 499394
rect 66322 499158 102086 499394
rect 102322 499158 138086 499394
rect 138322 499158 174086 499394
rect 174322 499158 210086 499394
rect 210322 499158 246086 499394
rect 246322 499158 282086 499394
rect 282322 499158 318086 499394
rect 318322 499158 354086 499394
rect 354322 499158 390086 499394
rect 390322 499158 426086 499394
rect 426322 499158 462086 499394
rect 462322 499158 498086 499394
rect 498322 499158 534086 499394
rect 534322 499158 570086 499394
rect 570322 499158 592062 499394
rect 592298 499158 592382 499394
rect 592618 499158 592650 499394
rect -8726 498976 592650 499158
rect -6806 495694 590730 495876
rect -6806 495458 -6774 495694
rect -6538 495458 -6454 495694
rect -6218 495458 26386 495694
rect 26622 495458 62386 495694
rect 62622 495458 98386 495694
rect 98622 495458 134386 495694
rect 134622 495458 170386 495694
rect 170622 495458 206386 495694
rect 206622 495458 242386 495694
rect 242622 495458 278386 495694
rect 278622 495458 314386 495694
rect 314622 495458 350386 495694
rect 350622 495458 386386 495694
rect 386622 495458 422386 495694
rect 422622 495458 458386 495694
rect 458622 495458 494386 495694
rect 494622 495458 530386 495694
rect 530622 495458 566386 495694
rect 566622 495458 590142 495694
rect 590378 495458 590462 495694
rect 590698 495458 590730 495694
rect -6806 495276 590730 495458
rect -4886 491994 588810 492176
rect -4886 491758 -4854 491994
rect -4618 491758 -4534 491994
rect -4298 491758 22686 491994
rect 22922 491758 58686 491994
rect 58922 491758 94686 491994
rect 94922 491758 130686 491994
rect 130922 491758 166686 491994
rect 166922 491758 202686 491994
rect 202922 491758 238686 491994
rect 238922 491758 274686 491994
rect 274922 491758 310686 491994
rect 310922 491758 346686 491994
rect 346922 491758 382686 491994
rect 382922 491758 418686 491994
rect 418922 491758 454686 491994
rect 454922 491758 490686 491994
rect 490922 491758 526686 491994
rect 526922 491758 562686 491994
rect 562922 491758 588222 491994
rect 588458 491758 588542 491994
rect 588778 491758 588810 491994
rect -4886 491576 588810 491758
rect -2966 488294 586890 488476
rect -2966 488058 -2934 488294
rect -2698 488058 -2614 488294
rect -2378 488058 18986 488294
rect 19222 488058 54986 488294
rect 55222 488058 90986 488294
rect 91222 488058 126986 488294
rect 127222 488058 162986 488294
rect 163222 488058 198986 488294
rect 199222 488058 234986 488294
rect 235222 488058 270986 488294
rect 271222 488058 306986 488294
rect 307222 488058 342986 488294
rect 343222 488058 378986 488294
rect 379222 488058 414986 488294
rect 415222 488058 450986 488294
rect 451222 488058 486986 488294
rect 487222 488058 522986 488294
rect 523222 488058 558986 488294
rect 559222 488058 586302 488294
rect 586538 488058 586622 488294
rect 586858 488058 586890 488294
rect -2966 487876 586890 488058
rect -8726 481394 592650 481576
rect -8726 481158 -7734 481394
rect -7498 481158 -7414 481394
rect -7178 481158 12086 481394
rect 12322 481158 48086 481394
rect 48322 481158 84086 481394
rect 84322 481158 120086 481394
rect 120322 481158 156086 481394
rect 156322 481158 192086 481394
rect 192322 481158 228086 481394
rect 228322 481158 264086 481394
rect 264322 481158 300086 481394
rect 300322 481158 336086 481394
rect 336322 481158 372086 481394
rect 372322 481158 408086 481394
rect 408322 481158 444086 481394
rect 444322 481158 480086 481394
rect 480322 481158 516086 481394
rect 516322 481158 552086 481394
rect 552322 481158 591102 481394
rect 591338 481158 591422 481394
rect 591658 481158 592650 481394
rect -8726 480976 592650 481158
rect -6806 477694 590730 477876
rect -6806 477458 -5814 477694
rect -5578 477458 -5494 477694
rect -5258 477458 8386 477694
rect 8622 477458 44386 477694
rect 44622 477458 80386 477694
rect 80622 477458 116386 477694
rect 116622 477458 152386 477694
rect 152622 477458 188386 477694
rect 188622 477458 224386 477694
rect 224622 477458 260386 477694
rect 260622 477458 296386 477694
rect 296622 477458 332386 477694
rect 332622 477458 368386 477694
rect 368622 477458 404386 477694
rect 404622 477458 440386 477694
rect 440622 477458 476386 477694
rect 476622 477458 512386 477694
rect 512622 477458 548386 477694
rect 548622 477458 589182 477694
rect 589418 477458 589502 477694
rect 589738 477458 590730 477694
rect -6806 477276 590730 477458
rect -4886 473994 588810 474176
rect -4886 473758 -3894 473994
rect -3658 473758 -3574 473994
rect -3338 473758 4686 473994
rect 4922 473758 40686 473994
rect 40922 473758 76686 473994
rect 76922 473758 112686 473994
rect 112922 473758 148686 473994
rect 148922 473758 184686 473994
rect 184922 473758 220686 473994
rect 220922 473758 256686 473994
rect 256922 473758 292686 473994
rect 292922 473758 328686 473994
rect 328922 473758 364686 473994
rect 364922 473758 400686 473994
rect 400922 473758 436686 473994
rect 436922 473758 472686 473994
rect 472922 473758 508686 473994
rect 508922 473758 544686 473994
rect 544922 473758 580686 473994
rect 580922 473758 587262 473994
rect 587498 473758 587582 473994
rect 587818 473758 588810 473994
rect -4886 473576 588810 473758
rect -2966 470294 586890 470476
rect -2966 470058 -1974 470294
rect -1738 470058 -1654 470294
rect -1418 470058 986 470294
rect 1222 470058 36986 470294
rect 37222 470058 72986 470294
rect 73222 470058 108986 470294
rect 109222 470058 144986 470294
rect 145222 470058 180986 470294
rect 181222 470058 216986 470294
rect 217222 470058 252986 470294
rect 253222 470058 288986 470294
rect 289222 470058 324986 470294
rect 325222 470058 360986 470294
rect 361222 470058 396986 470294
rect 397222 470058 432986 470294
rect 433222 470058 468986 470294
rect 469222 470058 504986 470294
rect 505222 470058 540986 470294
rect 541222 470058 576986 470294
rect 577222 470058 585342 470294
rect 585578 470058 585662 470294
rect 585898 470058 586890 470294
rect -2966 469876 586890 470058
rect -8726 463394 592650 463576
rect -8726 463158 -8694 463394
rect -8458 463158 -8374 463394
rect -8138 463158 30086 463394
rect 30322 463158 66086 463394
rect 66322 463158 102086 463394
rect 102322 463158 138086 463394
rect 138322 463158 174086 463394
rect 174322 463158 210086 463394
rect 210322 463158 246086 463394
rect 246322 463158 282086 463394
rect 282322 463158 318086 463394
rect 318322 463158 354086 463394
rect 354322 463158 390086 463394
rect 390322 463158 426086 463394
rect 426322 463158 462086 463394
rect 462322 463158 498086 463394
rect 498322 463158 534086 463394
rect 534322 463158 570086 463394
rect 570322 463158 592062 463394
rect 592298 463158 592382 463394
rect 592618 463158 592650 463394
rect -8726 462976 592650 463158
rect -6806 459694 590730 459876
rect -6806 459458 -6774 459694
rect -6538 459458 -6454 459694
rect -6218 459458 26386 459694
rect 26622 459458 62386 459694
rect 62622 459458 98386 459694
rect 98622 459458 134386 459694
rect 134622 459458 170386 459694
rect 170622 459458 206386 459694
rect 206622 459458 242386 459694
rect 242622 459458 278386 459694
rect 278622 459458 314386 459694
rect 314622 459458 350386 459694
rect 350622 459458 386386 459694
rect 386622 459458 422386 459694
rect 422622 459458 458386 459694
rect 458622 459458 494386 459694
rect 494622 459458 530386 459694
rect 530622 459458 566386 459694
rect 566622 459458 590142 459694
rect 590378 459458 590462 459694
rect 590698 459458 590730 459694
rect -6806 459276 590730 459458
rect -4886 455994 588810 456176
rect -4886 455758 -4854 455994
rect -4618 455758 -4534 455994
rect -4298 455758 22686 455994
rect 22922 455758 58686 455994
rect 58922 455758 94686 455994
rect 94922 455758 130686 455994
rect 130922 455758 166686 455994
rect 166922 455758 202686 455994
rect 202922 455758 238686 455994
rect 238922 455758 274686 455994
rect 274922 455758 310686 455994
rect 310922 455758 346686 455994
rect 346922 455758 382686 455994
rect 382922 455758 418686 455994
rect 418922 455758 454686 455994
rect 454922 455758 490686 455994
rect 490922 455758 526686 455994
rect 526922 455758 562686 455994
rect 562922 455758 588222 455994
rect 588458 455758 588542 455994
rect 588778 455758 588810 455994
rect -4886 455576 588810 455758
rect -2966 452294 586890 452476
rect -2966 452058 -2934 452294
rect -2698 452058 -2614 452294
rect -2378 452058 18986 452294
rect 19222 452058 54986 452294
rect 55222 452058 90986 452294
rect 91222 452058 126986 452294
rect 127222 452058 162986 452294
rect 163222 452058 198986 452294
rect 199222 452058 234986 452294
rect 235222 452058 270986 452294
rect 271222 452058 306986 452294
rect 307222 452058 342986 452294
rect 343222 452058 378986 452294
rect 379222 452058 414986 452294
rect 415222 452058 450986 452294
rect 451222 452058 486986 452294
rect 487222 452058 522986 452294
rect 523222 452058 558986 452294
rect 559222 452058 586302 452294
rect 586538 452058 586622 452294
rect 586858 452058 586890 452294
rect -2966 451876 586890 452058
rect -8726 445394 592650 445576
rect -8726 445158 -7734 445394
rect -7498 445158 -7414 445394
rect -7178 445158 12086 445394
rect 12322 445158 48086 445394
rect 48322 445158 84086 445394
rect 84322 445158 120086 445394
rect 120322 445158 156086 445394
rect 156322 445158 192086 445394
rect 192322 445158 228086 445394
rect 228322 445158 264086 445394
rect 264322 445158 300086 445394
rect 300322 445158 336086 445394
rect 336322 445158 372086 445394
rect 372322 445158 408086 445394
rect 408322 445158 444086 445394
rect 444322 445158 480086 445394
rect 480322 445158 516086 445394
rect 516322 445158 552086 445394
rect 552322 445158 591102 445394
rect 591338 445158 591422 445394
rect 591658 445158 592650 445394
rect -8726 444976 592650 445158
rect -6806 441694 590730 441876
rect -6806 441458 -5814 441694
rect -5578 441458 -5494 441694
rect -5258 441458 8386 441694
rect 8622 441458 44386 441694
rect 44622 441458 80386 441694
rect 80622 441458 116386 441694
rect 116622 441458 152386 441694
rect 152622 441458 188386 441694
rect 188622 441458 224386 441694
rect 224622 441458 260386 441694
rect 260622 441458 296386 441694
rect 296622 441458 332386 441694
rect 332622 441458 368386 441694
rect 368622 441458 404386 441694
rect 404622 441458 440386 441694
rect 440622 441458 476386 441694
rect 476622 441458 512386 441694
rect 512622 441458 548386 441694
rect 548622 441458 589182 441694
rect 589418 441458 589502 441694
rect 589738 441458 590730 441694
rect -6806 441276 590730 441458
rect -4886 437994 588810 438176
rect -4886 437758 -3894 437994
rect -3658 437758 -3574 437994
rect -3338 437758 4686 437994
rect 4922 437758 40686 437994
rect 40922 437758 76686 437994
rect 76922 437758 112686 437994
rect 112922 437758 148686 437994
rect 148922 437758 184686 437994
rect 184922 437758 220686 437994
rect 220922 437758 256686 437994
rect 256922 437758 292686 437994
rect 292922 437758 328686 437994
rect 328922 437758 364686 437994
rect 364922 437758 400686 437994
rect 400922 437758 436686 437994
rect 436922 437758 472686 437994
rect 472922 437758 508686 437994
rect 508922 437758 544686 437994
rect 544922 437758 580686 437994
rect 580922 437758 587262 437994
rect 587498 437758 587582 437994
rect 587818 437758 588810 437994
rect -4886 437576 588810 437758
rect -2966 434294 586890 434476
rect -2966 434058 -1974 434294
rect -1738 434058 -1654 434294
rect -1418 434058 986 434294
rect 1222 434058 36986 434294
rect 37222 434058 72986 434294
rect 73222 434058 108986 434294
rect 109222 434058 144986 434294
rect 145222 434058 180986 434294
rect 181222 434058 216986 434294
rect 217222 434058 252986 434294
rect 253222 434058 288986 434294
rect 289222 434058 324986 434294
rect 325222 434058 360986 434294
rect 361222 434058 396986 434294
rect 397222 434058 432986 434294
rect 433222 434058 468986 434294
rect 469222 434058 504986 434294
rect 505222 434058 540986 434294
rect 541222 434058 576986 434294
rect 577222 434058 585342 434294
rect 585578 434058 585662 434294
rect 585898 434058 586890 434294
rect -2966 433876 586890 434058
rect -8726 427394 592650 427576
rect -8726 427158 -8694 427394
rect -8458 427158 -8374 427394
rect -8138 427158 30086 427394
rect 30322 427158 66086 427394
rect 66322 427158 102086 427394
rect 102322 427158 138086 427394
rect 138322 427158 174086 427394
rect 174322 427158 210086 427394
rect 210322 427158 246086 427394
rect 246322 427158 282086 427394
rect 282322 427158 318086 427394
rect 318322 427158 354086 427394
rect 354322 427158 390086 427394
rect 390322 427158 426086 427394
rect 426322 427158 462086 427394
rect 462322 427158 498086 427394
rect 498322 427158 534086 427394
rect 534322 427158 570086 427394
rect 570322 427158 592062 427394
rect 592298 427158 592382 427394
rect 592618 427158 592650 427394
rect -8726 426976 592650 427158
rect -6806 423694 590730 423876
rect -6806 423458 -6774 423694
rect -6538 423458 -6454 423694
rect -6218 423458 26386 423694
rect 26622 423458 206386 423694
rect 206622 423458 242386 423694
rect 242622 423458 278386 423694
rect 278622 423458 314386 423694
rect 314622 423458 494386 423694
rect 494622 423458 530386 423694
rect 530622 423458 566386 423694
rect 566622 423458 590142 423694
rect 590378 423458 590462 423694
rect 590698 423458 590730 423694
rect -6806 423276 590730 423458
rect -4886 419994 588810 420176
rect -4886 419758 -4854 419994
rect -4618 419758 -4534 419994
rect -4298 419758 22686 419994
rect 22922 419758 202686 419994
rect 202922 419758 238686 419994
rect 238922 419758 274686 419994
rect 274922 419758 310686 419994
rect 310922 419758 490686 419994
rect 490922 419758 526686 419994
rect 526922 419758 562686 419994
rect 562922 419758 588222 419994
rect 588458 419758 588542 419994
rect 588778 419758 588810 419994
rect -4886 419576 588810 419758
rect -2966 416294 586890 416476
rect -2966 416058 -2934 416294
rect -2698 416058 -2614 416294
rect -2378 416058 18986 416294
rect 19222 416058 40328 416294
rect 40564 416058 176056 416294
rect 176292 416058 198986 416294
rect 199222 416058 234986 416294
rect 235222 416058 270986 416294
rect 271222 416058 306986 416294
rect 307222 416058 340328 416294
rect 340564 416058 476056 416294
rect 476292 416058 486986 416294
rect 487222 416058 522986 416294
rect 523222 416058 558986 416294
rect 559222 416058 586302 416294
rect 586538 416058 586622 416294
rect 586858 416058 586890 416294
rect -2966 415876 586890 416058
rect -8726 409394 592650 409576
rect -8726 409158 -7734 409394
rect -7498 409158 -7414 409394
rect -7178 409158 12086 409394
rect 12322 409158 192086 409394
rect 192322 409158 228086 409394
rect 228322 409158 264086 409394
rect 264322 409158 300086 409394
rect 300322 409158 336086 409394
rect 336322 409158 480086 409394
rect 480322 409158 516086 409394
rect 516322 409158 552086 409394
rect 552322 409158 591102 409394
rect 591338 409158 591422 409394
rect 591658 409158 592650 409394
rect -8726 408976 592650 409158
rect -6806 405694 590730 405876
rect -6806 405458 -5814 405694
rect -5578 405458 -5494 405694
rect -5258 405458 8386 405694
rect 8622 405458 188386 405694
rect 188622 405458 224386 405694
rect 224622 405458 260386 405694
rect 260622 405458 296386 405694
rect 296622 405458 332386 405694
rect 332622 405458 512386 405694
rect 512622 405458 548386 405694
rect 548622 405458 589182 405694
rect 589418 405458 589502 405694
rect 589738 405458 590730 405694
rect -6806 405276 590730 405458
rect -4886 401994 588810 402176
rect -4886 401758 -3894 401994
rect -3658 401758 -3574 401994
rect -3338 401758 4686 401994
rect 4922 401758 184686 401994
rect 184922 401758 220686 401994
rect 220922 401758 256686 401994
rect 256922 401758 292686 401994
rect 292922 401758 328686 401994
rect 328922 401758 508686 401994
rect 508922 401758 544686 401994
rect 544922 401758 580686 401994
rect 580922 401758 587262 401994
rect 587498 401758 587582 401994
rect 587818 401758 588810 401994
rect -4886 401576 588810 401758
rect -2966 398294 586890 398476
rect -2966 398058 -1974 398294
rect -1738 398058 -1654 398294
rect -1418 398058 986 398294
rect 1222 398058 36986 398294
rect 37222 398058 41008 398294
rect 41244 398058 175376 398294
rect 175612 398058 180986 398294
rect 181222 398058 216986 398294
rect 217222 398058 252986 398294
rect 253222 398058 288986 398294
rect 289222 398058 324986 398294
rect 325222 398058 341008 398294
rect 341244 398058 475376 398294
rect 475612 398058 504986 398294
rect 505222 398058 540986 398294
rect 541222 398058 576986 398294
rect 577222 398058 585342 398294
rect 585578 398058 585662 398294
rect 585898 398058 586890 398294
rect -2966 397876 586890 398058
rect -8726 391394 592650 391576
rect -8726 391158 -8694 391394
rect -8458 391158 -8374 391394
rect -8138 391158 30086 391394
rect 30322 391158 210086 391394
rect 210322 391158 246086 391394
rect 246322 391158 282086 391394
rect 282322 391158 318086 391394
rect 318322 391158 498086 391394
rect 498322 391158 534086 391394
rect 534322 391158 570086 391394
rect 570322 391158 592062 391394
rect 592298 391158 592382 391394
rect 592618 391158 592650 391394
rect -8726 390976 592650 391158
rect -6806 387694 590730 387876
rect -6806 387458 -6774 387694
rect -6538 387458 -6454 387694
rect -6218 387458 26386 387694
rect 26622 387458 206386 387694
rect 206622 387458 242386 387694
rect 242622 387458 278386 387694
rect 278622 387458 314386 387694
rect 314622 387458 494386 387694
rect 494622 387458 530386 387694
rect 530622 387458 566386 387694
rect 566622 387458 590142 387694
rect 590378 387458 590462 387694
rect 590698 387458 590730 387694
rect -6806 387276 590730 387458
rect -4886 383994 588810 384176
rect -4886 383758 -4854 383994
rect -4618 383758 -4534 383994
rect -4298 383758 22686 383994
rect 22922 383758 202686 383994
rect 202922 383758 238686 383994
rect 238922 383758 274686 383994
rect 274922 383758 310686 383994
rect 310922 383758 490686 383994
rect 490922 383758 526686 383994
rect 526922 383758 562686 383994
rect 562922 383758 588222 383994
rect 588458 383758 588542 383994
rect 588778 383758 588810 383994
rect -4886 383576 588810 383758
rect -2966 380294 586890 380476
rect -2966 380058 -2934 380294
rect -2698 380058 -2614 380294
rect -2378 380058 18986 380294
rect 19222 380058 40328 380294
rect 40564 380058 176056 380294
rect 176292 380058 198986 380294
rect 199222 380058 234986 380294
rect 235222 380058 270986 380294
rect 271222 380058 306986 380294
rect 307222 380058 340328 380294
rect 340564 380058 476056 380294
rect 476292 380058 486986 380294
rect 487222 380058 522986 380294
rect 523222 380058 558986 380294
rect 559222 380058 586302 380294
rect 586538 380058 586622 380294
rect 586858 380058 586890 380294
rect -2966 379876 586890 380058
rect -8726 373394 592650 373576
rect -8726 373158 -7734 373394
rect -7498 373158 -7414 373394
rect -7178 373158 12086 373394
rect 12322 373158 192086 373394
rect 192322 373158 228086 373394
rect 228322 373158 264086 373394
rect 264322 373158 300086 373394
rect 300322 373158 336086 373394
rect 336322 373158 480086 373394
rect 480322 373158 516086 373394
rect 516322 373158 552086 373394
rect 552322 373158 591102 373394
rect 591338 373158 591422 373394
rect 591658 373158 592650 373394
rect -8726 372976 592650 373158
rect -6806 369694 590730 369876
rect -6806 369458 -5814 369694
rect -5578 369458 -5494 369694
rect -5258 369458 8386 369694
rect 8622 369458 188386 369694
rect 188622 369458 224386 369694
rect 224622 369458 260386 369694
rect 260622 369458 296386 369694
rect 296622 369458 332386 369694
rect 332622 369458 512386 369694
rect 512622 369458 548386 369694
rect 548622 369458 589182 369694
rect 589418 369458 589502 369694
rect 589738 369458 590730 369694
rect -6806 369276 590730 369458
rect -4886 365994 588810 366176
rect -4886 365758 -3894 365994
rect -3658 365758 -3574 365994
rect -3338 365758 4686 365994
rect 4922 365758 184686 365994
rect 184922 365758 220686 365994
rect 220922 365758 256686 365994
rect 256922 365758 292686 365994
rect 292922 365758 328686 365994
rect 328922 365758 508686 365994
rect 508922 365758 544686 365994
rect 544922 365758 580686 365994
rect 580922 365758 587262 365994
rect 587498 365758 587582 365994
rect 587818 365758 588810 365994
rect -4886 365576 588810 365758
rect -2966 362294 586890 362476
rect -2966 362058 -1974 362294
rect -1738 362058 -1654 362294
rect -1418 362058 986 362294
rect 1222 362058 36986 362294
rect 37222 362058 41008 362294
rect 41244 362058 175376 362294
rect 175612 362058 180986 362294
rect 181222 362058 216986 362294
rect 217222 362058 252986 362294
rect 253222 362058 288986 362294
rect 289222 362058 324986 362294
rect 325222 362058 341008 362294
rect 341244 362058 475376 362294
rect 475612 362058 504986 362294
rect 505222 362058 540986 362294
rect 541222 362058 576986 362294
rect 577222 362058 585342 362294
rect 585578 362058 585662 362294
rect 585898 362058 586890 362294
rect -2966 361876 586890 362058
rect -8726 355394 592650 355576
rect -8726 355158 -8694 355394
rect -8458 355158 -8374 355394
rect -8138 355158 30086 355394
rect 30322 355158 210086 355394
rect 210322 355158 246086 355394
rect 246322 355158 282086 355394
rect 282322 355158 318086 355394
rect 318322 355158 498086 355394
rect 498322 355158 534086 355394
rect 534322 355158 570086 355394
rect 570322 355158 592062 355394
rect 592298 355158 592382 355394
rect 592618 355158 592650 355394
rect -8726 354976 592650 355158
rect -6806 351694 590730 351876
rect -6806 351458 -6774 351694
rect -6538 351458 -6454 351694
rect -6218 351458 26386 351694
rect 26622 351458 206386 351694
rect 206622 351458 242386 351694
rect 242622 351458 278386 351694
rect 278622 351458 314386 351694
rect 314622 351458 494386 351694
rect 494622 351458 530386 351694
rect 530622 351458 566386 351694
rect 566622 351458 590142 351694
rect 590378 351458 590462 351694
rect 590698 351458 590730 351694
rect -6806 351276 590730 351458
rect -4886 347994 588810 348176
rect -4886 347758 -4854 347994
rect -4618 347758 -4534 347994
rect -4298 347758 22686 347994
rect 22922 347758 202686 347994
rect 202922 347758 238686 347994
rect 238922 347758 274686 347994
rect 274922 347758 310686 347994
rect 310922 347758 490686 347994
rect 490922 347758 526686 347994
rect 526922 347758 562686 347994
rect 562922 347758 588222 347994
rect 588458 347758 588542 347994
rect 588778 347758 588810 347994
rect -4886 347576 588810 347758
rect -2966 344294 586890 344476
rect -2966 344058 -2934 344294
rect -2698 344058 -2614 344294
rect -2378 344058 18986 344294
rect 19222 344058 40328 344294
rect 40564 344058 176056 344294
rect 176292 344058 198986 344294
rect 199222 344058 234986 344294
rect 235222 344058 270986 344294
rect 271222 344058 306986 344294
rect 307222 344058 340328 344294
rect 340564 344058 476056 344294
rect 476292 344058 486986 344294
rect 487222 344058 522986 344294
rect 523222 344058 558986 344294
rect 559222 344058 586302 344294
rect 586538 344058 586622 344294
rect 586858 344058 586890 344294
rect -2966 343876 586890 344058
rect -8726 337394 592650 337576
rect -8726 337158 -7734 337394
rect -7498 337158 -7414 337394
rect -7178 337158 12086 337394
rect 12322 337158 48086 337394
rect 48322 337158 84086 337394
rect 84322 337158 120086 337394
rect 120322 337158 156086 337394
rect 156322 337158 192086 337394
rect 192322 337158 228086 337394
rect 228322 337158 264086 337394
rect 264322 337158 300086 337394
rect 300322 337158 336086 337394
rect 336322 337158 372086 337394
rect 372322 337158 408086 337394
rect 408322 337158 444086 337394
rect 444322 337158 480086 337394
rect 480322 337158 516086 337394
rect 516322 337158 552086 337394
rect 552322 337158 591102 337394
rect 591338 337158 591422 337394
rect 591658 337158 592650 337394
rect -8726 336976 592650 337158
rect -6806 333694 590730 333876
rect -6806 333458 -5814 333694
rect -5578 333458 -5494 333694
rect -5258 333458 8386 333694
rect 8622 333458 44386 333694
rect 44622 333458 80386 333694
rect 80622 333458 116386 333694
rect 116622 333458 152386 333694
rect 152622 333458 188386 333694
rect 188622 333458 224386 333694
rect 224622 333458 260386 333694
rect 260622 333458 296386 333694
rect 296622 333458 332386 333694
rect 332622 333458 368386 333694
rect 368622 333458 404386 333694
rect 404622 333458 440386 333694
rect 440622 333458 476386 333694
rect 476622 333458 512386 333694
rect 512622 333458 548386 333694
rect 548622 333458 589182 333694
rect 589418 333458 589502 333694
rect 589738 333458 590730 333694
rect -6806 333276 590730 333458
rect -4886 329994 588810 330176
rect -4886 329758 -3894 329994
rect -3658 329758 -3574 329994
rect -3338 329758 4686 329994
rect 4922 329758 40686 329994
rect 40922 329758 76686 329994
rect 76922 329758 112686 329994
rect 112922 329758 148686 329994
rect 148922 329758 184686 329994
rect 184922 329758 220686 329994
rect 220922 329758 256686 329994
rect 256922 329758 292686 329994
rect 292922 329758 328686 329994
rect 328922 329758 364686 329994
rect 364922 329758 400686 329994
rect 400922 329758 436686 329994
rect 436922 329758 472686 329994
rect 472922 329758 508686 329994
rect 508922 329758 544686 329994
rect 544922 329758 580686 329994
rect 580922 329758 587262 329994
rect 587498 329758 587582 329994
rect 587818 329758 588810 329994
rect -4886 329576 588810 329758
rect -2966 326294 586890 326476
rect -2966 326058 -1974 326294
rect -1738 326058 -1654 326294
rect -1418 326058 986 326294
rect 1222 326058 36986 326294
rect 37222 326058 72986 326294
rect 73222 326058 108986 326294
rect 109222 326058 144986 326294
rect 145222 326058 180986 326294
rect 181222 326058 216986 326294
rect 217222 326058 252986 326294
rect 253222 326058 288986 326294
rect 289222 326058 324986 326294
rect 325222 326058 360986 326294
rect 361222 326058 396986 326294
rect 397222 326058 432986 326294
rect 433222 326058 468986 326294
rect 469222 326058 504986 326294
rect 505222 326058 540986 326294
rect 541222 326058 576986 326294
rect 577222 326058 585342 326294
rect 585578 326058 585662 326294
rect 585898 326058 586890 326294
rect -2966 325876 586890 326058
rect -8726 319394 592650 319576
rect -8726 319158 -8694 319394
rect -8458 319158 -8374 319394
rect -8138 319158 30086 319394
rect 30322 319158 66086 319394
rect 66322 319158 102086 319394
rect 102322 319158 138086 319394
rect 138322 319158 174086 319394
rect 174322 319158 210086 319394
rect 210322 319158 246086 319394
rect 246322 319158 282086 319394
rect 282322 319158 318086 319394
rect 318322 319158 354086 319394
rect 354322 319158 390086 319394
rect 390322 319158 426086 319394
rect 426322 319158 462086 319394
rect 462322 319158 498086 319394
rect 498322 319158 534086 319394
rect 534322 319158 570086 319394
rect 570322 319158 592062 319394
rect 592298 319158 592382 319394
rect 592618 319158 592650 319394
rect -8726 318976 592650 319158
rect -6806 315694 590730 315876
rect -6806 315458 -6774 315694
rect -6538 315458 -6454 315694
rect -6218 315458 26386 315694
rect 26622 315458 62386 315694
rect 62622 315458 98386 315694
rect 98622 315458 134386 315694
rect 134622 315458 170386 315694
rect 170622 315458 206386 315694
rect 206622 315458 242386 315694
rect 242622 315458 278386 315694
rect 278622 315458 314386 315694
rect 314622 315458 350386 315694
rect 350622 315458 386386 315694
rect 386622 315458 422386 315694
rect 422622 315458 458386 315694
rect 458622 315458 494386 315694
rect 494622 315458 530386 315694
rect 530622 315458 566386 315694
rect 566622 315458 590142 315694
rect 590378 315458 590462 315694
rect 590698 315458 590730 315694
rect -6806 315276 590730 315458
rect -4886 311994 588810 312176
rect -4886 311758 -4854 311994
rect -4618 311758 -4534 311994
rect -4298 311758 22686 311994
rect 22922 311758 58686 311994
rect 58922 311758 94686 311994
rect 94922 311758 130686 311994
rect 130922 311758 166686 311994
rect 166922 311758 202686 311994
rect 202922 311758 238686 311994
rect 238922 311758 274686 311994
rect 274922 311758 310686 311994
rect 310922 311758 346686 311994
rect 346922 311758 382686 311994
rect 382922 311758 418686 311994
rect 418922 311758 454686 311994
rect 454922 311758 490686 311994
rect 490922 311758 526686 311994
rect 526922 311758 562686 311994
rect 562922 311758 588222 311994
rect 588458 311758 588542 311994
rect 588778 311758 588810 311994
rect -4886 311576 588810 311758
rect -2966 308294 586890 308476
rect -2966 308058 -2934 308294
rect -2698 308058 -2614 308294
rect -2378 308058 18986 308294
rect 19222 308058 54986 308294
rect 55222 308058 90986 308294
rect 91222 308058 126986 308294
rect 127222 308058 162986 308294
rect 163222 308058 198986 308294
rect 199222 308058 234986 308294
rect 235222 308058 270986 308294
rect 271222 308058 306986 308294
rect 307222 308058 342986 308294
rect 343222 308058 378986 308294
rect 379222 308058 414986 308294
rect 415222 308058 450986 308294
rect 451222 308058 486986 308294
rect 487222 308058 522986 308294
rect 523222 308058 558986 308294
rect 559222 308058 586302 308294
rect 586538 308058 586622 308294
rect 586858 308058 586890 308294
rect -2966 307876 586890 308058
rect -8726 301394 592650 301576
rect -8726 301158 -7734 301394
rect -7498 301158 -7414 301394
rect -7178 301158 12086 301394
rect 12322 301158 48086 301394
rect 48322 301158 84086 301394
rect 84322 301158 120086 301394
rect 120322 301158 156086 301394
rect 156322 301158 192086 301394
rect 192322 301158 228086 301394
rect 228322 301158 264086 301394
rect 264322 301158 300086 301394
rect 300322 301158 336086 301394
rect 336322 301158 372086 301394
rect 372322 301158 408086 301394
rect 408322 301158 444086 301394
rect 444322 301158 480086 301394
rect 480322 301158 516086 301394
rect 516322 301158 552086 301394
rect 552322 301158 591102 301394
rect 591338 301158 591422 301394
rect 591658 301158 592650 301394
rect -8726 300976 592650 301158
rect -6806 297694 590730 297876
rect -6806 297458 -5814 297694
rect -5578 297458 -5494 297694
rect -5258 297458 8386 297694
rect 8622 297458 44386 297694
rect 44622 297458 80386 297694
rect 80622 297458 116386 297694
rect 116622 297458 152386 297694
rect 152622 297458 188386 297694
rect 188622 297458 224386 297694
rect 224622 297458 260386 297694
rect 260622 297458 296386 297694
rect 296622 297458 332386 297694
rect 332622 297458 368386 297694
rect 368622 297458 404386 297694
rect 404622 297458 440386 297694
rect 440622 297458 476386 297694
rect 476622 297458 512386 297694
rect 512622 297458 548386 297694
rect 548622 297458 589182 297694
rect 589418 297458 589502 297694
rect 589738 297458 590730 297694
rect -6806 297276 590730 297458
rect -4886 293994 588810 294176
rect -4886 293758 -3894 293994
rect -3658 293758 -3574 293994
rect -3338 293758 4686 293994
rect 4922 293758 40686 293994
rect 40922 293758 76686 293994
rect 76922 293758 112686 293994
rect 112922 293758 148686 293994
rect 148922 293758 184686 293994
rect 184922 293758 220686 293994
rect 220922 293758 256686 293994
rect 256922 293758 292686 293994
rect 292922 293758 328686 293994
rect 328922 293758 364686 293994
rect 364922 293758 400686 293994
rect 400922 293758 436686 293994
rect 436922 293758 472686 293994
rect 472922 293758 508686 293994
rect 508922 293758 544686 293994
rect 544922 293758 580686 293994
rect 580922 293758 587262 293994
rect 587498 293758 587582 293994
rect 587818 293758 588810 293994
rect -4886 293576 588810 293758
rect -2966 290294 586890 290476
rect -2966 290058 -1974 290294
rect -1738 290058 -1654 290294
rect -1418 290058 986 290294
rect 1222 290058 36986 290294
rect 37222 290058 72986 290294
rect 73222 290058 108986 290294
rect 109222 290058 144986 290294
rect 145222 290058 180986 290294
rect 181222 290058 216986 290294
rect 217222 290058 252986 290294
rect 253222 290058 288986 290294
rect 289222 290058 324986 290294
rect 325222 290058 360986 290294
rect 361222 290058 396986 290294
rect 397222 290058 432986 290294
rect 433222 290058 468986 290294
rect 469222 290058 504986 290294
rect 505222 290058 540986 290294
rect 541222 290058 576986 290294
rect 577222 290058 585342 290294
rect 585578 290058 585662 290294
rect 585898 290058 586890 290294
rect -2966 289876 586890 290058
rect -8726 283394 592650 283576
rect -8726 283158 -8694 283394
rect -8458 283158 -8374 283394
rect -8138 283158 30086 283394
rect 30322 283158 66086 283394
rect 66322 283158 102086 283394
rect 102322 283158 138086 283394
rect 138322 283158 174086 283394
rect 174322 283158 210086 283394
rect 210322 283158 246086 283394
rect 246322 283158 282086 283394
rect 282322 283158 318086 283394
rect 318322 283158 354086 283394
rect 354322 283158 390086 283394
rect 390322 283158 426086 283394
rect 426322 283158 462086 283394
rect 462322 283158 498086 283394
rect 498322 283158 534086 283394
rect 534322 283158 570086 283394
rect 570322 283158 592062 283394
rect 592298 283158 592382 283394
rect 592618 283158 592650 283394
rect -8726 282976 592650 283158
rect -6806 279694 590730 279876
rect -6806 279458 -6774 279694
rect -6538 279458 -6454 279694
rect -6218 279458 26386 279694
rect 26622 279458 62386 279694
rect 62622 279458 98386 279694
rect 98622 279458 134386 279694
rect 134622 279458 170386 279694
rect 170622 279458 206386 279694
rect 206622 279458 242386 279694
rect 242622 279458 278386 279694
rect 278622 279458 314386 279694
rect 314622 279458 350386 279694
rect 350622 279458 386386 279694
rect 386622 279458 422386 279694
rect 422622 279458 458386 279694
rect 458622 279458 494386 279694
rect 494622 279458 530386 279694
rect 530622 279458 566386 279694
rect 566622 279458 590142 279694
rect 590378 279458 590462 279694
rect 590698 279458 590730 279694
rect -6806 279276 590730 279458
rect -4886 275994 588810 276176
rect -4886 275758 -4854 275994
rect -4618 275758 -4534 275994
rect -4298 275758 22686 275994
rect 22922 275758 58686 275994
rect 58922 275758 94686 275994
rect 94922 275758 130686 275994
rect 130922 275758 166686 275994
rect 166922 275758 202686 275994
rect 202922 275758 238686 275994
rect 238922 275758 274686 275994
rect 274922 275758 310686 275994
rect 310922 275758 346686 275994
rect 346922 275758 382686 275994
rect 382922 275758 418686 275994
rect 418922 275758 454686 275994
rect 454922 275758 490686 275994
rect 490922 275758 526686 275994
rect 526922 275758 562686 275994
rect 562922 275758 588222 275994
rect 588458 275758 588542 275994
rect 588778 275758 588810 275994
rect -4886 275576 588810 275758
rect -2966 272294 586890 272476
rect -2966 272058 -2934 272294
rect -2698 272058 -2614 272294
rect -2378 272058 18986 272294
rect 19222 272058 54986 272294
rect 55222 272058 90986 272294
rect 91222 272058 126986 272294
rect 127222 272058 162986 272294
rect 163222 272058 198986 272294
rect 199222 272058 234986 272294
rect 235222 272058 270986 272294
rect 271222 272058 306986 272294
rect 307222 272058 342986 272294
rect 343222 272058 378986 272294
rect 379222 272058 414986 272294
rect 415222 272058 450986 272294
rect 451222 272058 486986 272294
rect 487222 272058 522986 272294
rect 523222 272058 558986 272294
rect 559222 272058 586302 272294
rect 586538 272058 586622 272294
rect 586858 272058 586890 272294
rect -2966 271876 586890 272058
rect -8726 265394 592650 265576
rect -8726 265158 -7734 265394
rect -7498 265158 -7414 265394
rect -7178 265158 12086 265394
rect 12322 265158 48086 265394
rect 48322 265158 84086 265394
rect 84322 265158 120086 265394
rect 120322 265158 156086 265394
rect 156322 265158 192086 265394
rect 192322 265158 228086 265394
rect 228322 265158 264086 265394
rect 264322 265158 300086 265394
rect 300322 265158 336086 265394
rect 336322 265158 372086 265394
rect 372322 265158 408086 265394
rect 408322 265158 444086 265394
rect 444322 265158 480086 265394
rect 480322 265158 516086 265394
rect 516322 265158 552086 265394
rect 552322 265158 591102 265394
rect 591338 265158 591422 265394
rect 591658 265158 592650 265394
rect -8726 264976 592650 265158
rect -6806 261694 590730 261876
rect -6806 261458 -5814 261694
rect -5578 261458 -5494 261694
rect -5258 261458 8386 261694
rect 8622 261458 44386 261694
rect 44622 261458 80386 261694
rect 80622 261458 116386 261694
rect 116622 261458 152386 261694
rect 152622 261458 188386 261694
rect 188622 261458 224386 261694
rect 224622 261458 260386 261694
rect 260622 261458 296386 261694
rect 296622 261458 332386 261694
rect 332622 261458 368386 261694
rect 368622 261458 404386 261694
rect 404622 261458 440386 261694
rect 440622 261458 476386 261694
rect 476622 261458 512386 261694
rect 512622 261458 548386 261694
rect 548622 261458 589182 261694
rect 589418 261458 589502 261694
rect 589738 261458 590730 261694
rect -6806 261276 590730 261458
rect -4886 257994 588810 258176
rect -4886 257758 -3894 257994
rect -3658 257758 -3574 257994
rect -3338 257758 4686 257994
rect 4922 257758 40686 257994
rect 40922 257758 76686 257994
rect 76922 257758 112686 257994
rect 112922 257758 148686 257994
rect 148922 257758 184686 257994
rect 184922 257758 220686 257994
rect 220922 257758 256686 257994
rect 256922 257758 292686 257994
rect 292922 257758 328686 257994
rect 328922 257758 364686 257994
rect 364922 257758 400686 257994
rect 400922 257758 436686 257994
rect 436922 257758 472686 257994
rect 472922 257758 508686 257994
rect 508922 257758 544686 257994
rect 544922 257758 580686 257994
rect 580922 257758 587262 257994
rect 587498 257758 587582 257994
rect 587818 257758 588810 257994
rect -4886 257576 588810 257758
rect -2966 254294 586890 254476
rect -2966 254058 -1974 254294
rect -1738 254058 -1654 254294
rect -1418 254058 986 254294
rect 1222 254058 36986 254294
rect 37222 254058 72986 254294
rect 73222 254058 108986 254294
rect 109222 254058 144986 254294
rect 145222 254058 180986 254294
rect 181222 254058 216986 254294
rect 217222 254058 252986 254294
rect 253222 254058 288986 254294
rect 289222 254058 324986 254294
rect 325222 254058 360986 254294
rect 361222 254058 396986 254294
rect 397222 254058 432986 254294
rect 433222 254058 468986 254294
rect 469222 254058 504986 254294
rect 505222 254058 540986 254294
rect 541222 254058 576986 254294
rect 577222 254058 585342 254294
rect 585578 254058 585662 254294
rect 585898 254058 586890 254294
rect -2966 253876 586890 254058
rect -8726 247394 592650 247576
rect -8726 247158 -8694 247394
rect -8458 247158 -8374 247394
rect -8138 247158 30086 247394
rect 30322 247158 66086 247394
rect 66322 247158 102086 247394
rect 102322 247158 138086 247394
rect 138322 247158 174086 247394
rect 174322 247158 210086 247394
rect 210322 247158 246086 247394
rect 246322 247158 282086 247394
rect 282322 247158 318086 247394
rect 318322 247158 354086 247394
rect 354322 247158 390086 247394
rect 390322 247158 426086 247394
rect 426322 247158 462086 247394
rect 462322 247158 498086 247394
rect 498322 247158 534086 247394
rect 534322 247158 570086 247394
rect 570322 247158 592062 247394
rect 592298 247158 592382 247394
rect 592618 247158 592650 247394
rect -8726 246976 592650 247158
rect -6806 243694 590730 243876
rect -6806 243458 -6774 243694
rect -6538 243458 -6454 243694
rect -6218 243458 26386 243694
rect 26622 243458 62386 243694
rect 62622 243458 98386 243694
rect 98622 243458 134386 243694
rect 134622 243458 170386 243694
rect 170622 243458 206386 243694
rect 206622 243458 242386 243694
rect 242622 243458 278386 243694
rect 278622 243458 314386 243694
rect 314622 243458 350386 243694
rect 350622 243458 386386 243694
rect 386622 243458 422386 243694
rect 422622 243458 458386 243694
rect 458622 243458 494386 243694
rect 494622 243458 530386 243694
rect 530622 243458 566386 243694
rect 566622 243458 590142 243694
rect 590378 243458 590462 243694
rect 590698 243458 590730 243694
rect -6806 243276 590730 243458
rect -4886 239994 588810 240176
rect -4886 239758 -4854 239994
rect -4618 239758 -4534 239994
rect -4298 239758 22686 239994
rect 22922 239758 274686 239994
rect 274922 239758 310686 239994
rect 310922 239758 346686 239994
rect 346922 239758 382686 239994
rect 382922 239758 418686 239994
rect 418922 239758 454686 239994
rect 454922 239758 490686 239994
rect 490922 239758 526686 239994
rect 526922 239758 562686 239994
rect 562922 239758 588222 239994
rect 588458 239758 588542 239994
rect 588778 239758 588810 239994
rect -4886 239576 588810 239758
rect -2966 236294 586890 236476
rect -2966 236058 -2934 236294
rect -2698 236058 -2614 236294
rect -2378 236058 18986 236294
rect 19222 236058 59610 236294
rect 59846 236058 90330 236294
rect 90566 236058 121050 236294
rect 121286 236058 151770 236294
rect 152006 236058 182490 236294
rect 182726 236058 213210 236294
rect 213446 236058 270986 236294
rect 271222 236058 306986 236294
rect 307222 236058 342986 236294
rect 343222 236058 378986 236294
rect 379222 236058 414986 236294
rect 415222 236058 450986 236294
rect 451222 236058 486986 236294
rect 487222 236058 522986 236294
rect 523222 236058 558986 236294
rect 559222 236058 586302 236294
rect 586538 236058 586622 236294
rect 586858 236058 586890 236294
rect -2966 235876 586890 236058
rect -8726 229394 592650 229576
rect -8726 229158 -7734 229394
rect -7498 229158 -7414 229394
rect -7178 229158 12086 229394
rect 12322 229158 264086 229394
rect 264322 229158 300086 229394
rect 300322 229158 336086 229394
rect 336322 229158 372086 229394
rect 372322 229158 408086 229394
rect 408322 229158 444086 229394
rect 444322 229158 480086 229394
rect 480322 229158 516086 229394
rect 516322 229158 552086 229394
rect 552322 229158 591102 229394
rect 591338 229158 591422 229394
rect 591658 229158 592650 229394
rect -8726 228976 592650 229158
rect -6806 225694 590730 225876
rect -6806 225458 -5814 225694
rect -5578 225458 -5494 225694
rect -5258 225458 8386 225694
rect 8622 225458 260386 225694
rect 260622 225458 296386 225694
rect 296622 225458 332386 225694
rect 332622 225458 368386 225694
rect 368622 225458 404386 225694
rect 404622 225458 440386 225694
rect 440622 225458 476386 225694
rect 476622 225458 512386 225694
rect 512622 225458 548386 225694
rect 548622 225458 589182 225694
rect 589418 225458 589502 225694
rect 589738 225458 590730 225694
rect -6806 225276 590730 225458
rect -4886 221994 588810 222176
rect -4886 221758 -3894 221994
rect -3658 221758 -3574 221994
rect -3338 221758 4686 221994
rect 4922 221758 256686 221994
rect 256922 221758 292686 221994
rect 292922 221758 328686 221994
rect 328922 221758 364686 221994
rect 364922 221758 400686 221994
rect 400922 221758 436686 221994
rect 436922 221758 472686 221994
rect 472922 221758 508686 221994
rect 508922 221758 544686 221994
rect 544922 221758 580686 221994
rect 580922 221758 587262 221994
rect 587498 221758 587582 221994
rect 587818 221758 588810 221994
rect -4886 221576 588810 221758
rect -2966 218294 586890 218476
rect -2966 218058 -1974 218294
rect -1738 218058 -1654 218294
rect -1418 218058 986 218294
rect 1222 218058 36986 218294
rect 37222 218058 44250 218294
rect 44486 218058 74970 218294
rect 75206 218058 105690 218294
rect 105926 218058 136410 218294
rect 136646 218058 167130 218294
rect 167366 218058 197850 218294
rect 198086 218058 228570 218294
rect 228806 218058 252986 218294
rect 253222 218058 288986 218294
rect 289222 218058 324986 218294
rect 325222 218058 360986 218294
rect 361222 218058 396986 218294
rect 397222 218058 432986 218294
rect 433222 218058 468986 218294
rect 469222 218058 504986 218294
rect 505222 218058 540986 218294
rect 541222 218058 576986 218294
rect 577222 218058 585342 218294
rect 585578 218058 585662 218294
rect 585898 218058 586890 218294
rect -2966 217876 586890 218058
rect -8726 211394 592650 211576
rect -8726 211158 -8694 211394
rect -8458 211158 -8374 211394
rect -8138 211158 30086 211394
rect 30322 211158 246086 211394
rect 246322 211158 282086 211394
rect 282322 211158 318086 211394
rect 318322 211158 354086 211394
rect 354322 211158 390086 211394
rect 390322 211158 426086 211394
rect 426322 211158 462086 211394
rect 462322 211158 498086 211394
rect 498322 211158 534086 211394
rect 534322 211158 570086 211394
rect 570322 211158 592062 211394
rect 592298 211158 592382 211394
rect 592618 211158 592650 211394
rect -8726 210976 592650 211158
rect -6806 207694 590730 207876
rect -6806 207458 -6774 207694
rect -6538 207458 -6454 207694
rect -6218 207458 26386 207694
rect 26622 207458 242386 207694
rect 242622 207458 278386 207694
rect 278622 207458 314386 207694
rect 314622 207458 350386 207694
rect 350622 207458 386386 207694
rect 386622 207458 422386 207694
rect 422622 207458 458386 207694
rect 458622 207458 494386 207694
rect 494622 207458 530386 207694
rect 530622 207458 566386 207694
rect 566622 207458 590142 207694
rect 590378 207458 590462 207694
rect 590698 207458 590730 207694
rect -6806 207276 590730 207458
rect -4886 203994 588810 204176
rect -4886 203758 -4854 203994
rect -4618 203758 -4534 203994
rect -4298 203758 22686 203994
rect 22922 203758 274686 203994
rect 274922 203758 310686 203994
rect 310922 203758 346686 203994
rect 346922 203758 382686 203994
rect 382922 203758 418686 203994
rect 418922 203758 454686 203994
rect 454922 203758 490686 203994
rect 490922 203758 526686 203994
rect 526922 203758 562686 203994
rect 562922 203758 588222 203994
rect 588458 203758 588542 203994
rect 588778 203758 588810 203994
rect -4886 203576 588810 203758
rect -2966 200294 586890 200476
rect -2966 200058 -2934 200294
rect -2698 200058 -2614 200294
rect -2378 200058 18986 200294
rect 19222 200058 59610 200294
rect 59846 200058 90330 200294
rect 90566 200058 121050 200294
rect 121286 200058 151770 200294
rect 152006 200058 182490 200294
rect 182726 200058 213210 200294
rect 213446 200058 270986 200294
rect 271222 200058 306986 200294
rect 307222 200058 342986 200294
rect 343222 200058 378986 200294
rect 379222 200058 414986 200294
rect 415222 200058 450986 200294
rect 451222 200058 486986 200294
rect 487222 200058 522986 200294
rect 523222 200058 558986 200294
rect 559222 200058 586302 200294
rect 586538 200058 586622 200294
rect 586858 200058 586890 200294
rect -2966 199876 586890 200058
rect -8726 193394 592650 193576
rect -8726 193158 -7734 193394
rect -7498 193158 -7414 193394
rect -7178 193158 12086 193394
rect 12322 193158 264086 193394
rect 264322 193158 300086 193394
rect 300322 193158 336086 193394
rect 336322 193158 372086 193394
rect 372322 193158 408086 193394
rect 408322 193158 444086 193394
rect 444322 193158 480086 193394
rect 480322 193158 516086 193394
rect 516322 193158 552086 193394
rect 552322 193158 591102 193394
rect 591338 193158 591422 193394
rect 591658 193158 592650 193394
rect -8726 192976 592650 193158
rect -6806 189694 590730 189876
rect -6806 189458 -5814 189694
rect -5578 189458 -5494 189694
rect -5258 189458 8386 189694
rect 8622 189458 260386 189694
rect 260622 189458 296386 189694
rect 296622 189458 332386 189694
rect 332622 189458 368386 189694
rect 368622 189458 404386 189694
rect 404622 189458 440386 189694
rect 440622 189458 476386 189694
rect 476622 189458 512386 189694
rect 512622 189458 548386 189694
rect 548622 189458 589182 189694
rect 589418 189458 589502 189694
rect 589738 189458 590730 189694
rect -6806 189276 590730 189458
rect -4886 185994 588810 186176
rect -4886 185758 -3894 185994
rect -3658 185758 -3574 185994
rect -3338 185758 4686 185994
rect 4922 185758 256686 185994
rect 256922 185758 292686 185994
rect 292922 185758 328686 185994
rect 328922 185758 364686 185994
rect 364922 185758 400686 185994
rect 400922 185758 436686 185994
rect 436922 185758 472686 185994
rect 472922 185758 508686 185994
rect 508922 185758 544686 185994
rect 544922 185758 580686 185994
rect 580922 185758 587262 185994
rect 587498 185758 587582 185994
rect 587818 185758 588810 185994
rect -4886 185576 588810 185758
rect -2966 182294 586890 182476
rect -2966 182058 -1974 182294
rect -1738 182058 -1654 182294
rect -1418 182058 986 182294
rect 1222 182058 36986 182294
rect 37222 182058 44250 182294
rect 44486 182058 74970 182294
rect 75206 182058 105690 182294
rect 105926 182058 136410 182294
rect 136646 182058 167130 182294
rect 167366 182058 197850 182294
rect 198086 182058 228570 182294
rect 228806 182058 252986 182294
rect 253222 182058 288986 182294
rect 289222 182058 324986 182294
rect 325222 182058 360986 182294
rect 361222 182058 396986 182294
rect 397222 182058 432986 182294
rect 433222 182058 468986 182294
rect 469222 182058 504986 182294
rect 505222 182058 540986 182294
rect 541222 182058 576986 182294
rect 577222 182058 585342 182294
rect 585578 182058 585662 182294
rect 585898 182058 586890 182294
rect -2966 181876 586890 182058
rect -8726 175394 592650 175576
rect -8726 175158 -8694 175394
rect -8458 175158 -8374 175394
rect -8138 175158 30086 175394
rect 30322 175158 246086 175394
rect 246322 175158 282086 175394
rect 282322 175158 318086 175394
rect 318322 175158 354086 175394
rect 354322 175158 390086 175394
rect 390322 175158 426086 175394
rect 426322 175158 462086 175394
rect 462322 175158 498086 175394
rect 498322 175158 534086 175394
rect 534322 175158 570086 175394
rect 570322 175158 592062 175394
rect 592298 175158 592382 175394
rect 592618 175158 592650 175394
rect -8726 174976 592650 175158
rect -6806 171694 590730 171876
rect -6806 171458 -6774 171694
rect -6538 171458 -6454 171694
rect -6218 171458 26386 171694
rect 26622 171458 242386 171694
rect 242622 171458 278386 171694
rect 278622 171458 314386 171694
rect 314622 171458 350386 171694
rect 350622 171458 386386 171694
rect 386622 171458 422386 171694
rect 422622 171458 458386 171694
rect 458622 171458 494386 171694
rect 494622 171458 530386 171694
rect 530622 171458 566386 171694
rect 566622 171458 590142 171694
rect 590378 171458 590462 171694
rect 590698 171458 590730 171694
rect -6806 171276 590730 171458
rect -4886 167994 588810 168176
rect -4886 167758 -4854 167994
rect -4618 167758 -4534 167994
rect -4298 167758 22686 167994
rect 22922 167758 274686 167994
rect 274922 167758 310686 167994
rect 310922 167758 346686 167994
rect 346922 167758 382686 167994
rect 382922 167758 418686 167994
rect 418922 167758 454686 167994
rect 454922 167758 490686 167994
rect 490922 167758 526686 167994
rect 526922 167758 562686 167994
rect 562922 167758 588222 167994
rect 588458 167758 588542 167994
rect 588778 167758 588810 167994
rect -4886 167576 588810 167758
rect -2966 164294 586890 164476
rect -2966 164058 -2934 164294
rect -2698 164058 -2614 164294
rect -2378 164058 18986 164294
rect 19222 164058 59610 164294
rect 59846 164058 90330 164294
rect 90566 164058 121050 164294
rect 121286 164058 151770 164294
rect 152006 164058 182490 164294
rect 182726 164058 213210 164294
rect 213446 164058 270986 164294
rect 271222 164058 306986 164294
rect 307222 164058 342986 164294
rect 343222 164058 378986 164294
rect 379222 164058 414986 164294
rect 415222 164058 450986 164294
rect 451222 164058 486986 164294
rect 487222 164058 522986 164294
rect 523222 164058 558986 164294
rect 559222 164058 586302 164294
rect 586538 164058 586622 164294
rect 586858 164058 586890 164294
rect -2966 163876 586890 164058
rect -8726 157394 592650 157576
rect -8726 157158 -7734 157394
rect -7498 157158 -7414 157394
rect -7178 157158 12086 157394
rect 12322 157158 264086 157394
rect 264322 157158 300086 157394
rect 300322 157158 336086 157394
rect 336322 157158 372086 157394
rect 372322 157158 408086 157394
rect 408322 157158 444086 157394
rect 444322 157158 480086 157394
rect 480322 157158 516086 157394
rect 516322 157158 552086 157394
rect 552322 157158 591102 157394
rect 591338 157158 591422 157394
rect 591658 157158 592650 157394
rect -8726 156976 592650 157158
rect -6806 153694 590730 153876
rect -6806 153458 -5814 153694
rect -5578 153458 -5494 153694
rect -5258 153458 8386 153694
rect 8622 153458 260386 153694
rect 260622 153458 296386 153694
rect 296622 153458 332386 153694
rect 332622 153458 368386 153694
rect 368622 153458 404386 153694
rect 404622 153458 440386 153694
rect 440622 153458 476386 153694
rect 476622 153458 512386 153694
rect 512622 153458 548386 153694
rect 548622 153458 589182 153694
rect 589418 153458 589502 153694
rect 589738 153458 590730 153694
rect -6806 153276 590730 153458
rect -4886 149994 588810 150176
rect -4886 149758 -3894 149994
rect -3658 149758 -3574 149994
rect -3338 149758 4686 149994
rect 4922 149758 256686 149994
rect 256922 149758 292686 149994
rect 292922 149758 328686 149994
rect 328922 149758 364686 149994
rect 364922 149758 400686 149994
rect 400922 149758 436686 149994
rect 436922 149758 472686 149994
rect 472922 149758 508686 149994
rect 508922 149758 544686 149994
rect 544922 149758 580686 149994
rect 580922 149758 587262 149994
rect 587498 149758 587582 149994
rect 587818 149758 588810 149994
rect -4886 149576 588810 149758
rect -2966 146294 586890 146476
rect -2966 146058 -1974 146294
rect -1738 146058 -1654 146294
rect -1418 146058 986 146294
rect 1222 146058 36986 146294
rect 37222 146058 44250 146294
rect 44486 146058 74970 146294
rect 75206 146058 105690 146294
rect 105926 146058 136410 146294
rect 136646 146058 167130 146294
rect 167366 146058 197850 146294
rect 198086 146058 228570 146294
rect 228806 146058 252986 146294
rect 253222 146058 288986 146294
rect 289222 146058 324986 146294
rect 325222 146058 360986 146294
rect 361222 146058 396986 146294
rect 397222 146058 432986 146294
rect 433222 146058 468986 146294
rect 469222 146058 504986 146294
rect 505222 146058 540986 146294
rect 541222 146058 576986 146294
rect 577222 146058 585342 146294
rect 585578 146058 585662 146294
rect 585898 146058 586890 146294
rect -2966 145876 586890 146058
rect -8726 139394 592650 139576
rect -8726 139158 -8694 139394
rect -8458 139158 -8374 139394
rect -8138 139158 30086 139394
rect 30322 139158 246086 139394
rect 246322 139158 282086 139394
rect 282322 139158 318086 139394
rect 318322 139158 354086 139394
rect 354322 139158 390086 139394
rect 390322 139158 426086 139394
rect 426322 139158 462086 139394
rect 462322 139158 498086 139394
rect 498322 139158 534086 139394
rect 534322 139158 570086 139394
rect 570322 139158 592062 139394
rect 592298 139158 592382 139394
rect 592618 139158 592650 139394
rect -8726 138976 592650 139158
rect -6806 135694 590730 135876
rect -6806 135458 -6774 135694
rect -6538 135458 -6454 135694
rect -6218 135458 26386 135694
rect 26622 135458 242386 135694
rect 242622 135458 278386 135694
rect 278622 135458 314386 135694
rect 314622 135458 350386 135694
rect 350622 135458 386386 135694
rect 386622 135458 422386 135694
rect 422622 135458 458386 135694
rect 458622 135458 494386 135694
rect 494622 135458 530386 135694
rect 530622 135458 566386 135694
rect 566622 135458 590142 135694
rect 590378 135458 590462 135694
rect 590698 135458 590730 135694
rect -6806 135276 590730 135458
rect -4886 131994 588810 132176
rect -4886 131758 -4854 131994
rect -4618 131758 -4534 131994
rect -4298 131758 22686 131994
rect 22922 131758 274686 131994
rect 274922 131758 310686 131994
rect 310922 131758 346686 131994
rect 346922 131758 382686 131994
rect 382922 131758 418686 131994
rect 418922 131758 454686 131994
rect 454922 131758 490686 131994
rect 490922 131758 526686 131994
rect 526922 131758 562686 131994
rect 562922 131758 588222 131994
rect 588458 131758 588542 131994
rect 588778 131758 588810 131994
rect -4886 131576 588810 131758
rect -2966 128294 586890 128476
rect -2966 128058 -2934 128294
rect -2698 128058 -2614 128294
rect -2378 128058 18986 128294
rect 19222 128058 59610 128294
rect 59846 128058 90330 128294
rect 90566 128058 121050 128294
rect 121286 128058 151770 128294
rect 152006 128058 182490 128294
rect 182726 128058 213210 128294
rect 213446 128058 270986 128294
rect 271222 128058 306986 128294
rect 307222 128058 342986 128294
rect 343222 128058 378986 128294
rect 379222 128058 414986 128294
rect 415222 128058 450986 128294
rect 451222 128058 486986 128294
rect 487222 128058 522986 128294
rect 523222 128058 558986 128294
rect 559222 128058 586302 128294
rect 586538 128058 586622 128294
rect 586858 128058 586890 128294
rect -2966 127876 586890 128058
rect -8726 121394 592650 121576
rect -8726 121158 -7734 121394
rect -7498 121158 -7414 121394
rect -7178 121158 12086 121394
rect 12322 121158 264086 121394
rect 264322 121158 300086 121394
rect 300322 121158 336086 121394
rect 336322 121158 372086 121394
rect 372322 121158 408086 121394
rect 408322 121158 444086 121394
rect 444322 121158 480086 121394
rect 480322 121158 516086 121394
rect 516322 121158 552086 121394
rect 552322 121158 591102 121394
rect 591338 121158 591422 121394
rect 591658 121158 592650 121394
rect -8726 120976 592650 121158
rect -6806 117694 590730 117876
rect -6806 117458 -5814 117694
rect -5578 117458 -5494 117694
rect -5258 117458 8386 117694
rect 8622 117458 260386 117694
rect 260622 117458 296386 117694
rect 296622 117458 332386 117694
rect 332622 117458 368386 117694
rect 368622 117458 404386 117694
rect 404622 117458 440386 117694
rect 440622 117458 476386 117694
rect 476622 117458 512386 117694
rect 512622 117458 548386 117694
rect 548622 117458 589182 117694
rect 589418 117458 589502 117694
rect 589738 117458 590730 117694
rect -6806 117276 590730 117458
rect -4886 113994 588810 114176
rect -4886 113758 -3894 113994
rect -3658 113758 -3574 113994
rect -3338 113758 4686 113994
rect 4922 113758 256686 113994
rect 256922 113758 292686 113994
rect 292922 113758 328686 113994
rect 328922 113758 364686 113994
rect 364922 113758 400686 113994
rect 400922 113758 436686 113994
rect 436922 113758 472686 113994
rect 472922 113758 508686 113994
rect 508922 113758 544686 113994
rect 544922 113758 580686 113994
rect 580922 113758 587262 113994
rect 587498 113758 587582 113994
rect 587818 113758 588810 113994
rect -4886 113576 588810 113758
rect -2966 110294 586890 110476
rect -2966 110058 -1974 110294
rect -1738 110058 -1654 110294
rect -1418 110058 986 110294
rect 1222 110058 36986 110294
rect 37222 110058 44250 110294
rect 44486 110058 74970 110294
rect 75206 110058 105690 110294
rect 105926 110058 136410 110294
rect 136646 110058 167130 110294
rect 167366 110058 197850 110294
rect 198086 110058 228570 110294
rect 228806 110058 252986 110294
rect 253222 110058 288986 110294
rect 289222 110058 324986 110294
rect 325222 110058 360986 110294
rect 361222 110058 396986 110294
rect 397222 110058 432986 110294
rect 433222 110058 468986 110294
rect 469222 110058 504986 110294
rect 505222 110058 540986 110294
rect 541222 110058 576986 110294
rect 577222 110058 585342 110294
rect 585578 110058 585662 110294
rect 585898 110058 586890 110294
rect -2966 109876 586890 110058
rect -8726 103394 592650 103576
rect -8726 103158 -8694 103394
rect -8458 103158 -8374 103394
rect -8138 103158 30086 103394
rect 30322 103158 246086 103394
rect 246322 103158 282086 103394
rect 282322 103158 318086 103394
rect 318322 103158 354086 103394
rect 354322 103158 390086 103394
rect 390322 103158 426086 103394
rect 426322 103158 462086 103394
rect 462322 103158 498086 103394
rect 498322 103158 534086 103394
rect 534322 103158 570086 103394
rect 570322 103158 592062 103394
rect 592298 103158 592382 103394
rect 592618 103158 592650 103394
rect -8726 102976 592650 103158
rect -6806 99694 590730 99876
rect -6806 99458 -6774 99694
rect -6538 99458 -6454 99694
rect -6218 99458 26386 99694
rect 26622 99458 242386 99694
rect 242622 99458 278386 99694
rect 278622 99458 314386 99694
rect 314622 99458 350386 99694
rect 350622 99458 386386 99694
rect 386622 99458 422386 99694
rect 422622 99458 458386 99694
rect 458622 99458 494386 99694
rect 494622 99458 530386 99694
rect 530622 99458 566386 99694
rect 566622 99458 590142 99694
rect 590378 99458 590462 99694
rect 590698 99458 590730 99694
rect -6806 99276 590730 99458
rect -4886 95994 588810 96176
rect -4886 95758 -4854 95994
rect -4618 95758 -4534 95994
rect -4298 95758 22686 95994
rect 22922 95758 274686 95994
rect 274922 95758 310686 95994
rect 310922 95758 346686 95994
rect 346922 95758 382686 95994
rect 382922 95758 418686 95994
rect 418922 95758 454686 95994
rect 454922 95758 490686 95994
rect 490922 95758 526686 95994
rect 526922 95758 562686 95994
rect 562922 95758 588222 95994
rect 588458 95758 588542 95994
rect 588778 95758 588810 95994
rect -4886 95576 588810 95758
rect -2966 92294 586890 92476
rect -2966 92058 -2934 92294
rect -2698 92058 -2614 92294
rect -2378 92058 18986 92294
rect 19222 92058 59610 92294
rect 59846 92058 90330 92294
rect 90566 92058 121050 92294
rect 121286 92058 151770 92294
rect 152006 92058 182490 92294
rect 182726 92058 213210 92294
rect 213446 92058 270986 92294
rect 271222 92058 306986 92294
rect 307222 92058 342986 92294
rect 343222 92058 378986 92294
rect 379222 92058 414986 92294
rect 415222 92058 450986 92294
rect 451222 92058 486986 92294
rect 487222 92058 522986 92294
rect 523222 92058 558986 92294
rect 559222 92058 586302 92294
rect 586538 92058 586622 92294
rect 586858 92058 586890 92294
rect -2966 91876 586890 92058
rect -8726 85394 592650 85576
rect -8726 85158 -7734 85394
rect -7498 85158 -7414 85394
rect -7178 85158 12086 85394
rect 12322 85158 264086 85394
rect 264322 85158 300086 85394
rect 300322 85158 336086 85394
rect 336322 85158 372086 85394
rect 372322 85158 408086 85394
rect 408322 85158 444086 85394
rect 444322 85158 480086 85394
rect 480322 85158 516086 85394
rect 516322 85158 552086 85394
rect 552322 85158 591102 85394
rect 591338 85158 591422 85394
rect 591658 85158 592650 85394
rect -8726 84976 592650 85158
rect -6806 81694 590730 81876
rect -6806 81458 -5814 81694
rect -5578 81458 -5494 81694
rect -5258 81458 8386 81694
rect 8622 81458 260386 81694
rect 260622 81458 296386 81694
rect 296622 81458 332386 81694
rect 332622 81458 368386 81694
rect 368622 81458 404386 81694
rect 404622 81458 440386 81694
rect 440622 81458 476386 81694
rect 476622 81458 512386 81694
rect 512622 81458 548386 81694
rect 548622 81458 589182 81694
rect 589418 81458 589502 81694
rect 589738 81458 590730 81694
rect -6806 81276 590730 81458
rect -4886 77994 588810 78176
rect -4886 77758 -3894 77994
rect -3658 77758 -3574 77994
rect -3338 77758 4686 77994
rect 4922 77758 256686 77994
rect 256922 77758 292686 77994
rect 292922 77758 328686 77994
rect 328922 77758 364686 77994
rect 364922 77758 400686 77994
rect 400922 77758 436686 77994
rect 436922 77758 472686 77994
rect 472922 77758 508686 77994
rect 508922 77758 544686 77994
rect 544922 77758 580686 77994
rect 580922 77758 587262 77994
rect 587498 77758 587582 77994
rect 587818 77758 588810 77994
rect -4886 77576 588810 77758
rect -2966 74294 586890 74476
rect -2966 74058 -1974 74294
rect -1738 74058 -1654 74294
rect -1418 74058 986 74294
rect 1222 74058 36986 74294
rect 37222 74058 44250 74294
rect 44486 74058 74970 74294
rect 75206 74058 105690 74294
rect 105926 74058 136410 74294
rect 136646 74058 167130 74294
rect 167366 74058 197850 74294
rect 198086 74058 228570 74294
rect 228806 74058 252986 74294
rect 253222 74058 288986 74294
rect 289222 74058 324986 74294
rect 325222 74058 360986 74294
rect 361222 74058 396986 74294
rect 397222 74058 432986 74294
rect 433222 74058 468986 74294
rect 469222 74058 504986 74294
rect 505222 74058 540986 74294
rect 541222 74058 576986 74294
rect 577222 74058 585342 74294
rect 585578 74058 585662 74294
rect 585898 74058 586890 74294
rect -2966 73876 586890 74058
rect -8726 67394 592650 67576
rect -8726 67158 -8694 67394
rect -8458 67158 -8374 67394
rect -8138 67158 30086 67394
rect 30322 67158 246086 67394
rect 246322 67158 282086 67394
rect 282322 67158 318086 67394
rect 318322 67158 354086 67394
rect 354322 67158 390086 67394
rect 390322 67158 426086 67394
rect 426322 67158 462086 67394
rect 462322 67158 498086 67394
rect 498322 67158 534086 67394
rect 534322 67158 570086 67394
rect 570322 67158 592062 67394
rect 592298 67158 592382 67394
rect 592618 67158 592650 67394
rect -8726 66976 592650 67158
rect -6806 63694 590730 63876
rect -6806 63458 -6774 63694
rect -6538 63458 -6454 63694
rect -6218 63458 26386 63694
rect 26622 63458 242386 63694
rect 242622 63458 278386 63694
rect 278622 63458 314386 63694
rect 314622 63458 350386 63694
rect 350622 63458 386386 63694
rect 386622 63458 422386 63694
rect 422622 63458 458386 63694
rect 458622 63458 494386 63694
rect 494622 63458 530386 63694
rect 530622 63458 566386 63694
rect 566622 63458 590142 63694
rect 590378 63458 590462 63694
rect 590698 63458 590730 63694
rect -6806 63276 590730 63458
rect -4886 59994 588810 60176
rect -4886 59758 -4854 59994
rect -4618 59758 -4534 59994
rect -4298 59758 22686 59994
rect 22922 59758 274686 59994
rect 274922 59758 310686 59994
rect 310922 59758 346686 59994
rect 346922 59758 382686 59994
rect 382922 59758 418686 59994
rect 418922 59758 454686 59994
rect 454922 59758 490686 59994
rect 490922 59758 526686 59994
rect 526922 59758 562686 59994
rect 562922 59758 588222 59994
rect 588458 59758 588542 59994
rect 588778 59758 588810 59994
rect -4886 59576 588810 59758
rect -2966 56294 586890 56476
rect -2966 56058 -2934 56294
rect -2698 56058 -2614 56294
rect -2378 56058 18986 56294
rect 19222 56058 59610 56294
rect 59846 56058 90330 56294
rect 90566 56058 121050 56294
rect 121286 56058 151770 56294
rect 152006 56058 182490 56294
rect 182726 56058 213210 56294
rect 213446 56058 270986 56294
rect 271222 56058 306986 56294
rect 307222 56058 342986 56294
rect 343222 56058 378986 56294
rect 379222 56058 414986 56294
rect 415222 56058 450986 56294
rect 451222 56058 486986 56294
rect 487222 56058 522986 56294
rect 523222 56058 558986 56294
rect 559222 56058 586302 56294
rect 586538 56058 586622 56294
rect 586858 56058 586890 56294
rect -2966 55876 586890 56058
rect -8726 49394 592650 49576
rect -8726 49158 -7734 49394
rect -7498 49158 -7414 49394
rect -7178 49158 12086 49394
rect 12322 49158 264086 49394
rect 264322 49158 300086 49394
rect 300322 49158 336086 49394
rect 336322 49158 372086 49394
rect 372322 49158 408086 49394
rect 408322 49158 444086 49394
rect 444322 49158 480086 49394
rect 480322 49158 516086 49394
rect 516322 49158 552086 49394
rect 552322 49158 591102 49394
rect 591338 49158 591422 49394
rect 591658 49158 592650 49394
rect -8726 48976 592650 49158
rect -6806 45694 590730 45876
rect -6806 45458 -5814 45694
rect -5578 45458 -5494 45694
rect -5258 45458 8386 45694
rect 8622 45458 260386 45694
rect 260622 45458 296386 45694
rect 296622 45458 332386 45694
rect 332622 45458 368386 45694
rect 368622 45458 404386 45694
rect 404622 45458 440386 45694
rect 440622 45458 476386 45694
rect 476622 45458 512386 45694
rect 512622 45458 548386 45694
rect 548622 45458 589182 45694
rect 589418 45458 589502 45694
rect 589738 45458 590730 45694
rect -6806 45276 590730 45458
rect -4886 41994 588810 42176
rect -4886 41758 -3894 41994
rect -3658 41758 -3574 41994
rect -3338 41758 4686 41994
rect 4922 41758 256686 41994
rect 256922 41758 292686 41994
rect 292922 41758 328686 41994
rect 328922 41758 364686 41994
rect 364922 41758 400686 41994
rect 400922 41758 436686 41994
rect 436922 41758 472686 41994
rect 472922 41758 508686 41994
rect 508922 41758 544686 41994
rect 544922 41758 580686 41994
rect 580922 41758 587262 41994
rect 587498 41758 587582 41994
rect 587818 41758 588810 41994
rect -4886 41576 588810 41758
rect -2966 38294 586890 38476
rect -2966 38058 -1974 38294
rect -1738 38058 -1654 38294
rect -1418 38058 986 38294
rect 1222 38058 36986 38294
rect 37222 38058 252986 38294
rect 253222 38058 288986 38294
rect 289222 38058 324986 38294
rect 325222 38058 360986 38294
rect 361222 38058 396986 38294
rect 397222 38058 432986 38294
rect 433222 38058 468986 38294
rect 469222 38058 504986 38294
rect 505222 38058 540986 38294
rect 541222 38058 576986 38294
rect 577222 38058 585342 38294
rect 585578 38058 585662 38294
rect 585898 38058 586890 38294
rect -2966 37876 586890 38058
rect -8726 31394 592650 31576
rect -8726 31158 -8694 31394
rect -8458 31158 -8374 31394
rect -8138 31158 30086 31394
rect 30322 31158 66086 31394
rect 66322 31158 102086 31394
rect 102322 31158 138086 31394
rect 138322 31158 174086 31394
rect 174322 31158 210086 31394
rect 210322 31158 246086 31394
rect 246322 31158 282086 31394
rect 282322 31158 318086 31394
rect 318322 31158 354086 31394
rect 354322 31158 390086 31394
rect 390322 31158 426086 31394
rect 426322 31158 462086 31394
rect 462322 31158 498086 31394
rect 498322 31158 534086 31394
rect 534322 31158 570086 31394
rect 570322 31158 592062 31394
rect 592298 31158 592382 31394
rect 592618 31158 592650 31394
rect -8726 30976 592650 31158
rect -6806 27694 590730 27876
rect -6806 27458 -6774 27694
rect -6538 27458 -6454 27694
rect -6218 27458 26386 27694
rect 26622 27458 62386 27694
rect 62622 27458 98386 27694
rect 98622 27458 134386 27694
rect 134622 27458 170386 27694
rect 170622 27458 206386 27694
rect 206622 27458 242386 27694
rect 242622 27458 278386 27694
rect 278622 27458 314386 27694
rect 314622 27458 350386 27694
rect 350622 27458 386386 27694
rect 386622 27458 422386 27694
rect 422622 27458 458386 27694
rect 458622 27458 494386 27694
rect 494622 27458 530386 27694
rect 530622 27458 566386 27694
rect 566622 27458 590142 27694
rect 590378 27458 590462 27694
rect 590698 27458 590730 27694
rect -6806 27276 590730 27458
rect -4886 23994 588810 24176
rect -4886 23758 -4854 23994
rect -4618 23758 -4534 23994
rect -4298 23758 22686 23994
rect 22922 23758 58686 23994
rect 58922 23758 94686 23994
rect 94922 23758 130686 23994
rect 130922 23758 166686 23994
rect 166922 23758 202686 23994
rect 202922 23758 238686 23994
rect 238922 23758 274686 23994
rect 274922 23758 310686 23994
rect 310922 23758 346686 23994
rect 346922 23758 382686 23994
rect 382922 23758 418686 23994
rect 418922 23758 454686 23994
rect 454922 23758 490686 23994
rect 490922 23758 526686 23994
rect 526922 23758 562686 23994
rect 562922 23758 588222 23994
rect 588458 23758 588542 23994
rect 588778 23758 588810 23994
rect -4886 23576 588810 23758
rect -2966 20294 586890 20476
rect -2966 20058 -2934 20294
rect -2698 20058 -2614 20294
rect -2378 20058 18986 20294
rect 19222 20058 54986 20294
rect 55222 20058 90986 20294
rect 91222 20058 126986 20294
rect 127222 20058 162986 20294
rect 163222 20058 198986 20294
rect 199222 20058 234986 20294
rect 235222 20058 270986 20294
rect 271222 20058 306986 20294
rect 307222 20058 342986 20294
rect 343222 20058 378986 20294
rect 379222 20058 414986 20294
rect 415222 20058 450986 20294
rect 451222 20058 486986 20294
rect 487222 20058 522986 20294
rect 523222 20058 558986 20294
rect 559222 20058 586302 20294
rect 586538 20058 586622 20294
rect 586858 20058 586890 20294
rect -2966 19876 586890 20058
rect -8726 13394 592650 13576
rect -8726 13158 -7734 13394
rect -7498 13158 -7414 13394
rect -7178 13158 12086 13394
rect 12322 13158 48086 13394
rect 48322 13158 84086 13394
rect 84322 13158 120086 13394
rect 120322 13158 156086 13394
rect 156322 13158 192086 13394
rect 192322 13158 228086 13394
rect 228322 13158 264086 13394
rect 264322 13158 300086 13394
rect 300322 13158 336086 13394
rect 336322 13158 372086 13394
rect 372322 13158 408086 13394
rect 408322 13158 444086 13394
rect 444322 13158 480086 13394
rect 480322 13158 516086 13394
rect 516322 13158 552086 13394
rect 552322 13158 591102 13394
rect 591338 13158 591422 13394
rect 591658 13158 592650 13394
rect -8726 12976 592650 13158
rect -6806 9694 590730 9876
rect -6806 9458 -5814 9694
rect -5578 9458 -5494 9694
rect -5258 9458 8386 9694
rect 8622 9458 44386 9694
rect 44622 9458 80386 9694
rect 80622 9458 116386 9694
rect 116622 9458 152386 9694
rect 152622 9458 188386 9694
rect 188622 9458 224386 9694
rect 224622 9458 260386 9694
rect 260622 9458 296386 9694
rect 296622 9458 332386 9694
rect 332622 9458 368386 9694
rect 368622 9458 404386 9694
rect 404622 9458 440386 9694
rect 440622 9458 476386 9694
rect 476622 9458 512386 9694
rect 512622 9458 548386 9694
rect 548622 9458 589182 9694
rect 589418 9458 589502 9694
rect 589738 9458 590730 9694
rect -6806 9276 590730 9458
rect -4886 5994 588810 6176
rect -4886 5758 -3894 5994
rect -3658 5758 -3574 5994
rect -3338 5758 4686 5994
rect 4922 5758 40686 5994
rect 40922 5758 76686 5994
rect 76922 5758 112686 5994
rect 112922 5758 148686 5994
rect 148922 5758 184686 5994
rect 184922 5758 220686 5994
rect 220922 5758 256686 5994
rect 256922 5758 292686 5994
rect 292922 5758 328686 5994
rect 328922 5758 364686 5994
rect 364922 5758 400686 5994
rect 400922 5758 436686 5994
rect 436922 5758 472686 5994
rect 472922 5758 508686 5994
rect 508922 5758 544686 5994
rect 544922 5758 580686 5994
rect 580922 5758 587262 5994
rect 587498 5758 587582 5994
rect 587818 5758 588810 5994
rect -4886 5576 588810 5758
rect -2966 2294 586890 2476
rect -2966 2058 -1974 2294
rect -1738 2058 -1654 2294
rect -1418 2058 986 2294
rect 1222 2058 36986 2294
rect 37222 2058 72986 2294
rect 73222 2058 108986 2294
rect 109222 2058 144986 2294
rect 145222 2058 180986 2294
rect 181222 2058 216986 2294
rect 217222 2058 252986 2294
rect 253222 2058 288986 2294
rect 289222 2058 324986 2294
rect 325222 2058 360986 2294
rect 361222 2058 396986 2294
rect 397222 2058 432986 2294
rect 433222 2058 468986 2294
rect 469222 2058 504986 2294
rect 505222 2058 540986 2294
rect 541222 2058 576986 2294
rect 577222 2058 585342 2294
rect 585578 2058 585662 2294
rect 585898 2058 586890 2294
rect -2966 1876 586890 2058
rect -2006 -346 585930 -314
rect -2006 -582 -1974 -346
rect -1738 -582 -1654 -346
rect -1418 -582 986 -346
rect 1222 -582 36986 -346
rect 37222 -582 72986 -346
rect 73222 -582 108986 -346
rect 109222 -582 144986 -346
rect 145222 -582 180986 -346
rect 181222 -582 216986 -346
rect 217222 -582 252986 -346
rect 253222 -582 288986 -346
rect 289222 -582 324986 -346
rect 325222 -582 360986 -346
rect 361222 -582 396986 -346
rect 397222 -582 432986 -346
rect 433222 -582 468986 -346
rect 469222 -582 504986 -346
rect 505222 -582 540986 -346
rect 541222 -582 576986 -346
rect 577222 -582 585342 -346
rect 585578 -582 585662 -346
rect 585898 -582 585930 -346
rect -2006 -666 585930 -582
rect -2006 -902 -1974 -666
rect -1738 -902 -1654 -666
rect -1418 -902 986 -666
rect 1222 -902 36986 -666
rect 37222 -902 72986 -666
rect 73222 -902 108986 -666
rect 109222 -902 144986 -666
rect 145222 -902 180986 -666
rect 181222 -902 216986 -666
rect 217222 -902 252986 -666
rect 253222 -902 288986 -666
rect 289222 -902 324986 -666
rect 325222 -902 360986 -666
rect 361222 -902 396986 -666
rect 397222 -902 432986 -666
rect 433222 -902 468986 -666
rect 469222 -902 504986 -666
rect 505222 -902 540986 -666
rect 541222 -902 576986 -666
rect 577222 -902 585342 -666
rect 585578 -902 585662 -666
rect 585898 -902 585930 -666
rect -2006 -934 585930 -902
rect -2966 -1306 586890 -1274
rect -2966 -1542 -2934 -1306
rect -2698 -1542 -2614 -1306
rect -2378 -1542 18986 -1306
rect 19222 -1542 54986 -1306
rect 55222 -1542 90986 -1306
rect 91222 -1542 126986 -1306
rect 127222 -1542 162986 -1306
rect 163222 -1542 198986 -1306
rect 199222 -1542 234986 -1306
rect 235222 -1542 270986 -1306
rect 271222 -1542 306986 -1306
rect 307222 -1542 342986 -1306
rect 343222 -1542 378986 -1306
rect 379222 -1542 414986 -1306
rect 415222 -1542 450986 -1306
rect 451222 -1542 486986 -1306
rect 487222 -1542 522986 -1306
rect 523222 -1542 558986 -1306
rect 559222 -1542 586302 -1306
rect 586538 -1542 586622 -1306
rect 586858 -1542 586890 -1306
rect -2966 -1626 586890 -1542
rect -2966 -1862 -2934 -1626
rect -2698 -1862 -2614 -1626
rect -2378 -1862 18986 -1626
rect 19222 -1862 54986 -1626
rect 55222 -1862 90986 -1626
rect 91222 -1862 126986 -1626
rect 127222 -1862 162986 -1626
rect 163222 -1862 198986 -1626
rect 199222 -1862 234986 -1626
rect 235222 -1862 270986 -1626
rect 271222 -1862 306986 -1626
rect 307222 -1862 342986 -1626
rect 343222 -1862 378986 -1626
rect 379222 -1862 414986 -1626
rect 415222 -1862 450986 -1626
rect 451222 -1862 486986 -1626
rect 487222 -1862 522986 -1626
rect 523222 -1862 558986 -1626
rect 559222 -1862 586302 -1626
rect 586538 -1862 586622 -1626
rect 586858 -1862 586890 -1626
rect -2966 -1894 586890 -1862
rect -3926 -2266 587850 -2234
rect -3926 -2502 -3894 -2266
rect -3658 -2502 -3574 -2266
rect -3338 -2502 4686 -2266
rect 4922 -2502 40686 -2266
rect 40922 -2502 76686 -2266
rect 76922 -2502 112686 -2266
rect 112922 -2502 148686 -2266
rect 148922 -2502 184686 -2266
rect 184922 -2502 220686 -2266
rect 220922 -2502 256686 -2266
rect 256922 -2502 292686 -2266
rect 292922 -2502 328686 -2266
rect 328922 -2502 364686 -2266
rect 364922 -2502 400686 -2266
rect 400922 -2502 436686 -2266
rect 436922 -2502 472686 -2266
rect 472922 -2502 508686 -2266
rect 508922 -2502 544686 -2266
rect 544922 -2502 580686 -2266
rect 580922 -2502 587262 -2266
rect 587498 -2502 587582 -2266
rect 587818 -2502 587850 -2266
rect -3926 -2586 587850 -2502
rect -3926 -2822 -3894 -2586
rect -3658 -2822 -3574 -2586
rect -3338 -2822 4686 -2586
rect 4922 -2822 40686 -2586
rect 40922 -2822 76686 -2586
rect 76922 -2822 112686 -2586
rect 112922 -2822 148686 -2586
rect 148922 -2822 184686 -2586
rect 184922 -2822 220686 -2586
rect 220922 -2822 256686 -2586
rect 256922 -2822 292686 -2586
rect 292922 -2822 328686 -2586
rect 328922 -2822 364686 -2586
rect 364922 -2822 400686 -2586
rect 400922 -2822 436686 -2586
rect 436922 -2822 472686 -2586
rect 472922 -2822 508686 -2586
rect 508922 -2822 544686 -2586
rect 544922 -2822 580686 -2586
rect 580922 -2822 587262 -2586
rect 587498 -2822 587582 -2586
rect 587818 -2822 587850 -2586
rect -3926 -2854 587850 -2822
rect -4886 -3226 588810 -3194
rect -4886 -3462 -4854 -3226
rect -4618 -3462 -4534 -3226
rect -4298 -3462 22686 -3226
rect 22922 -3462 58686 -3226
rect 58922 -3462 94686 -3226
rect 94922 -3462 130686 -3226
rect 130922 -3462 166686 -3226
rect 166922 -3462 202686 -3226
rect 202922 -3462 238686 -3226
rect 238922 -3462 274686 -3226
rect 274922 -3462 310686 -3226
rect 310922 -3462 346686 -3226
rect 346922 -3462 382686 -3226
rect 382922 -3462 418686 -3226
rect 418922 -3462 454686 -3226
rect 454922 -3462 490686 -3226
rect 490922 -3462 526686 -3226
rect 526922 -3462 562686 -3226
rect 562922 -3462 588222 -3226
rect 588458 -3462 588542 -3226
rect 588778 -3462 588810 -3226
rect -4886 -3546 588810 -3462
rect -4886 -3782 -4854 -3546
rect -4618 -3782 -4534 -3546
rect -4298 -3782 22686 -3546
rect 22922 -3782 58686 -3546
rect 58922 -3782 94686 -3546
rect 94922 -3782 130686 -3546
rect 130922 -3782 166686 -3546
rect 166922 -3782 202686 -3546
rect 202922 -3782 238686 -3546
rect 238922 -3782 274686 -3546
rect 274922 -3782 310686 -3546
rect 310922 -3782 346686 -3546
rect 346922 -3782 382686 -3546
rect 382922 -3782 418686 -3546
rect 418922 -3782 454686 -3546
rect 454922 -3782 490686 -3546
rect 490922 -3782 526686 -3546
rect 526922 -3782 562686 -3546
rect 562922 -3782 588222 -3546
rect 588458 -3782 588542 -3546
rect 588778 -3782 588810 -3546
rect -4886 -3814 588810 -3782
rect -5846 -4186 589770 -4154
rect -5846 -4422 -5814 -4186
rect -5578 -4422 -5494 -4186
rect -5258 -4422 8386 -4186
rect 8622 -4422 44386 -4186
rect 44622 -4422 80386 -4186
rect 80622 -4422 116386 -4186
rect 116622 -4422 152386 -4186
rect 152622 -4422 188386 -4186
rect 188622 -4422 224386 -4186
rect 224622 -4422 260386 -4186
rect 260622 -4422 296386 -4186
rect 296622 -4422 332386 -4186
rect 332622 -4422 368386 -4186
rect 368622 -4422 404386 -4186
rect 404622 -4422 440386 -4186
rect 440622 -4422 476386 -4186
rect 476622 -4422 512386 -4186
rect 512622 -4422 548386 -4186
rect 548622 -4422 589182 -4186
rect 589418 -4422 589502 -4186
rect 589738 -4422 589770 -4186
rect -5846 -4506 589770 -4422
rect -5846 -4742 -5814 -4506
rect -5578 -4742 -5494 -4506
rect -5258 -4742 8386 -4506
rect 8622 -4742 44386 -4506
rect 44622 -4742 80386 -4506
rect 80622 -4742 116386 -4506
rect 116622 -4742 152386 -4506
rect 152622 -4742 188386 -4506
rect 188622 -4742 224386 -4506
rect 224622 -4742 260386 -4506
rect 260622 -4742 296386 -4506
rect 296622 -4742 332386 -4506
rect 332622 -4742 368386 -4506
rect 368622 -4742 404386 -4506
rect 404622 -4742 440386 -4506
rect 440622 -4742 476386 -4506
rect 476622 -4742 512386 -4506
rect 512622 -4742 548386 -4506
rect 548622 -4742 589182 -4506
rect 589418 -4742 589502 -4506
rect 589738 -4742 589770 -4506
rect -5846 -4774 589770 -4742
rect -6806 -5146 590730 -5114
rect -6806 -5382 -6774 -5146
rect -6538 -5382 -6454 -5146
rect -6218 -5382 26386 -5146
rect 26622 -5382 62386 -5146
rect 62622 -5382 98386 -5146
rect 98622 -5382 134386 -5146
rect 134622 -5382 170386 -5146
rect 170622 -5382 206386 -5146
rect 206622 -5382 242386 -5146
rect 242622 -5382 278386 -5146
rect 278622 -5382 314386 -5146
rect 314622 -5382 350386 -5146
rect 350622 -5382 386386 -5146
rect 386622 -5382 422386 -5146
rect 422622 -5382 458386 -5146
rect 458622 -5382 494386 -5146
rect 494622 -5382 530386 -5146
rect 530622 -5382 566386 -5146
rect 566622 -5382 590142 -5146
rect 590378 -5382 590462 -5146
rect 590698 -5382 590730 -5146
rect -6806 -5466 590730 -5382
rect -6806 -5702 -6774 -5466
rect -6538 -5702 -6454 -5466
rect -6218 -5702 26386 -5466
rect 26622 -5702 62386 -5466
rect 62622 -5702 98386 -5466
rect 98622 -5702 134386 -5466
rect 134622 -5702 170386 -5466
rect 170622 -5702 206386 -5466
rect 206622 -5702 242386 -5466
rect 242622 -5702 278386 -5466
rect 278622 -5702 314386 -5466
rect 314622 -5702 350386 -5466
rect 350622 -5702 386386 -5466
rect 386622 -5702 422386 -5466
rect 422622 -5702 458386 -5466
rect 458622 -5702 494386 -5466
rect 494622 -5702 530386 -5466
rect 530622 -5702 566386 -5466
rect 566622 -5702 590142 -5466
rect 590378 -5702 590462 -5466
rect 590698 -5702 590730 -5466
rect -6806 -5734 590730 -5702
rect -7766 -6106 591690 -6074
rect -7766 -6342 -7734 -6106
rect -7498 -6342 -7414 -6106
rect -7178 -6342 12086 -6106
rect 12322 -6342 48086 -6106
rect 48322 -6342 84086 -6106
rect 84322 -6342 120086 -6106
rect 120322 -6342 156086 -6106
rect 156322 -6342 192086 -6106
rect 192322 -6342 228086 -6106
rect 228322 -6342 264086 -6106
rect 264322 -6342 300086 -6106
rect 300322 -6342 336086 -6106
rect 336322 -6342 372086 -6106
rect 372322 -6342 408086 -6106
rect 408322 -6342 444086 -6106
rect 444322 -6342 480086 -6106
rect 480322 -6342 516086 -6106
rect 516322 -6342 552086 -6106
rect 552322 -6342 591102 -6106
rect 591338 -6342 591422 -6106
rect 591658 -6342 591690 -6106
rect -7766 -6426 591690 -6342
rect -7766 -6662 -7734 -6426
rect -7498 -6662 -7414 -6426
rect -7178 -6662 12086 -6426
rect 12322 -6662 48086 -6426
rect 48322 -6662 84086 -6426
rect 84322 -6662 120086 -6426
rect 120322 -6662 156086 -6426
rect 156322 -6662 192086 -6426
rect 192322 -6662 228086 -6426
rect 228322 -6662 264086 -6426
rect 264322 -6662 300086 -6426
rect 300322 -6662 336086 -6426
rect 336322 -6662 372086 -6426
rect 372322 -6662 408086 -6426
rect 408322 -6662 444086 -6426
rect 444322 -6662 480086 -6426
rect 480322 -6662 516086 -6426
rect 516322 -6662 552086 -6426
rect 552322 -6662 591102 -6426
rect 591338 -6662 591422 -6426
rect 591658 -6662 591690 -6426
rect -7766 -6694 591690 -6662
rect -8726 -7066 592650 -7034
rect -8726 -7302 -8694 -7066
rect -8458 -7302 -8374 -7066
rect -8138 -7302 30086 -7066
rect 30322 -7302 66086 -7066
rect 66322 -7302 102086 -7066
rect 102322 -7302 138086 -7066
rect 138322 -7302 174086 -7066
rect 174322 -7302 210086 -7066
rect 210322 -7302 246086 -7066
rect 246322 -7302 282086 -7066
rect 282322 -7302 318086 -7066
rect 318322 -7302 354086 -7066
rect 354322 -7302 390086 -7066
rect 390322 -7302 426086 -7066
rect 426322 -7302 462086 -7066
rect 462322 -7302 498086 -7066
rect 498322 -7302 534086 -7066
rect 534322 -7302 570086 -7066
rect 570322 -7302 592062 -7066
rect 592298 -7302 592382 -7066
rect 592618 -7302 592650 -7066
rect -8726 -7386 592650 -7302
rect -8726 -7622 -8694 -7386
rect -8458 -7622 -8374 -7386
rect -8138 -7622 30086 -7386
rect 30322 -7622 66086 -7386
rect 66322 -7622 102086 -7386
rect 102322 -7622 138086 -7386
rect 138322 -7622 174086 -7386
rect 174322 -7622 210086 -7386
rect 210322 -7622 246086 -7386
rect 246322 -7622 282086 -7386
rect 282322 -7622 318086 -7386
rect 318322 -7622 354086 -7386
rect 354322 -7622 390086 -7386
rect 390322 -7622 426086 -7386
rect 426322 -7622 462086 -7386
rect 462322 -7622 498086 -7386
rect 498322 -7622 534086 -7386
rect 534322 -7622 570086 -7386
rect 570322 -7622 592062 -7386
rect 592298 -7622 592382 -7386
rect 592618 -7622 592650 -7386
rect -8726 -7654 592650 -7622
use sky130_sram_2kbyte_1rw1r_32x512_8  sram1
timestamp 1645332165
transform 1 0 340000 0 1 340000
box 0 0 136620 83308
use sky130_sram_2kbyte_1rw1r_32x512_8  sram
timestamp 1645332165
transform 1 0 40000 0 1 340000
box 0 0 136620 83308
use user_proj  mprj
timestamp 1645332165
transform 1 0 40000 0 1 40000
box 0 0 198160 200304
<< labels >>
rlabel metal3 s 583520 285276 584960 285516 6 analog_io[0]
port 0 nsew signal bidirectional
rlabel metal2 s 446098 703520 446210 704960 6 analog_io[10]
port 1 nsew signal bidirectional
rlabel metal2 s 381146 703520 381258 704960 6 analog_io[11]
port 2 nsew signal bidirectional
rlabel metal2 s 316286 703520 316398 704960 6 analog_io[12]
port 3 nsew signal bidirectional
rlabel metal2 s 251426 703520 251538 704960 6 analog_io[13]
port 4 nsew signal bidirectional
rlabel metal2 s 186474 703520 186586 704960 6 analog_io[14]
port 5 nsew signal bidirectional
rlabel metal2 s 121614 703520 121726 704960 6 analog_io[15]
port 6 nsew signal bidirectional
rlabel metal2 s 56754 703520 56866 704960 6 analog_io[16]
port 7 nsew signal bidirectional
rlabel metal3 s -960 697220 480 697460 4 analog_io[17]
port 8 nsew signal bidirectional
rlabel metal3 s -960 644996 480 645236 4 analog_io[18]
port 9 nsew signal bidirectional
rlabel metal3 s -960 592908 480 593148 4 analog_io[19]
port 10 nsew signal bidirectional
rlabel metal3 s 583520 338452 584960 338692 6 analog_io[1]
port 11 nsew signal bidirectional
rlabel metal3 s -960 540684 480 540924 4 analog_io[20]
port 12 nsew signal bidirectional
rlabel metal3 s -960 488596 480 488836 4 analog_io[21]
port 13 nsew signal bidirectional
rlabel metal3 s -960 436508 480 436748 4 analog_io[22]
port 14 nsew signal bidirectional
rlabel metal3 s -960 384284 480 384524 4 analog_io[23]
port 15 nsew signal bidirectional
rlabel metal3 s -960 332196 480 332436 4 analog_io[24]
port 16 nsew signal bidirectional
rlabel metal3 s -960 279972 480 280212 4 analog_io[25]
port 17 nsew signal bidirectional
rlabel metal3 s -960 227884 480 228124 4 analog_io[26]
port 18 nsew signal bidirectional
rlabel metal3 s -960 175796 480 176036 4 analog_io[27]
port 19 nsew signal bidirectional
rlabel metal3 s -960 123572 480 123812 4 analog_io[28]
port 20 nsew signal bidirectional
rlabel metal3 s 583520 391628 584960 391868 6 analog_io[2]
port 21 nsew signal bidirectional
rlabel metal3 s 583520 444668 584960 444908 6 analog_io[3]
port 22 nsew signal bidirectional
rlabel metal3 s 583520 497844 584960 498084 6 analog_io[4]
port 23 nsew signal bidirectional
rlabel metal3 s 583520 551020 584960 551260 6 analog_io[5]
port 24 nsew signal bidirectional
rlabel metal3 s 583520 604060 584960 604300 6 analog_io[6]
port 25 nsew signal bidirectional
rlabel metal3 s 583520 657236 584960 657476 6 analog_io[7]
port 26 nsew signal bidirectional
rlabel metal2 s 575818 703520 575930 704960 6 analog_io[8]
port 27 nsew signal bidirectional
rlabel metal2 s 510958 703520 511070 704960 6 analog_io[9]
port 28 nsew signal bidirectional
rlabel metal3 s 583520 6476 584960 6716 6 io_in[0]
port 29 nsew signal input
rlabel metal3 s 583520 457996 584960 458236 6 io_in[10]
port 30 nsew signal input
rlabel metal3 s 583520 511172 584960 511412 6 io_in[11]
port 31 nsew signal input
rlabel metal3 s 583520 564212 584960 564452 6 io_in[12]
port 32 nsew signal input
rlabel metal3 s 583520 617388 584960 617628 6 io_in[13]
port 33 nsew signal input
rlabel metal3 s 583520 670564 584960 670804 6 io_in[14]
port 34 nsew signal input
rlabel metal2 s 559626 703520 559738 704960 6 io_in[15]
port 35 nsew signal input
rlabel metal2 s 494766 703520 494878 704960 6 io_in[16]
port 36 nsew signal input
rlabel metal2 s 429814 703520 429926 704960 6 io_in[17]
port 37 nsew signal input
rlabel metal2 s 364954 703520 365066 704960 6 io_in[18]
port 38 nsew signal input
rlabel metal2 s 300094 703520 300206 704960 6 io_in[19]
port 39 nsew signal input
rlabel metal3 s 583520 46188 584960 46428 6 io_in[1]
port 40 nsew signal input
rlabel metal2 s 235142 703520 235254 704960 6 io_in[20]
port 41 nsew signal input
rlabel metal2 s 170282 703520 170394 704960 6 io_in[21]
port 42 nsew signal input
rlabel metal2 s 105422 703520 105534 704960 6 io_in[22]
port 43 nsew signal input
rlabel metal2 s 40470 703520 40582 704960 6 io_in[23]
port 44 nsew signal input
rlabel metal3 s -960 684164 480 684404 4 io_in[24]
port 45 nsew signal input
rlabel metal3 s -960 631940 480 632180 4 io_in[25]
port 46 nsew signal input
rlabel metal3 s -960 579852 480 580092 4 io_in[26]
port 47 nsew signal input
rlabel metal3 s -960 527764 480 528004 4 io_in[27]
port 48 nsew signal input
rlabel metal3 s -960 475540 480 475780 4 io_in[28]
port 49 nsew signal input
rlabel metal3 s -960 423452 480 423692 4 io_in[29]
port 50 nsew signal input
rlabel metal3 s 583520 86036 584960 86276 6 io_in[2]
port 51 nsew signal input
rlabel metal3 s -960 371228 480 371468 4 io_in[30]
port 52 nsew signal input
rlabel metal3 s -960 319140 480 319380 4 io_in[31]
port 53 nsew signal input
rlabel metal3 s -960 267052 480 267292 4 io_in[32]
port 54 nsew signal input
rlabel metal3 s -960 214828 480 215068 4 io_in[33]
port 55 nsew signal input
rlabel metal3 s -960 162740 480 162980 4 io_in[34]
port 56 nsew signal input
rlabel metal3 s -960 110516 480 110756 4 io_in[35]
port 57 nsew signal input
rlabel metal3 s -960 71484 480 71724 4 io_in[36]
port 58 nsew signal input
rlabel metal3 s -960 32316 480 32556 4 io_in[37]
port 59 nsew signal input
rlabel metal3 s 583520 125884 584960 126124 6 io_in[3]
port 60 nsew signal input
rlabel metal3 s 583520 165732 584960 165972 6 io_in[4]
port 61 nsew signal input
rlabel metal3 s 583520 205580 584960 205820 6 io_in[5]
port 62 nsew signal input
rlabel metal3 s 583520 245428 584960 245668 6 io_in[6]
port 63 nsew signal input
rlabel metal3 s 583520 298604 584960 298844 6 io_in[7]
port 64 nsew signal input
rlabel metal3 s 583520 351780 584960 352020 6 io_in[8]
port 65 nsew signal input
rlabel metal3 s 583520 404820 584960 405060 6 io_in[9]
port 66 nsew signal input
rlabel metal3 s 583520 32996 584960 33236 6 io_oeb[0]
port 67 nsew signal tristate
rlabel metal3 s 583520 484516 584960 484756 6 io_oeb[10]
port 68 nsew signal tristate
rlabel metal3 s 583520 537692 584960 537932 6 io_oeb[11]
port 69 nsew signal tristate
rlabel metal3 s 583520 590868 584960 591108 6 io_oeb[12]
port 70 nsew signal tristate
rlabel metal3 s 583520 643908 584960 644148 6 io_oeb[13]
port 71 nsew signal tristate
rlabel metal3 s 583520 697084 584960 697324 6 io_oeb[14]
port 72 nsew signal tristate
rlabel metal2 s 527150 703520 527262 704960 6 io_oeb[15]
port 73 nsew signal tristate
rlabel metal2 s 462290 703520 462402 704960 6 io_oeb[16]
port 74 nsew signal tristate
rlabel metal2 s 397430 703520 397542 704960 6 io_oeb[17]
port 75 nsew signal tristate
rlabel metal2 s 332478 703520 332590 704960 6 io_oeb[18]
port 76 nsew signal tristate
rlabel metal2 s 267618 703520 267730 704960 6 io_oeb[19]
port 77 nsew signal tristate
rlabel metal3 s 583520 72844 584960 73084 6 io_oeb[1]
port 78 nsew signal tristate
rlabel metal2 s 202758 703520 202870 704960 6 io_oeb[20]
port 79 nsew signal tristate
rlabel metal2 s 137806 703520 137918 704960 6 io_oeb[21]
port 80 nsew signal tristate
rlabel metal2 s 72946 703520 73058 704960 6 io_oeb[22]
port 81 nsew signal tristate
rlabel metal2 s 8086 703520 8198 704960 6 io_oeb[23]
port 82 nsew signal tristate
rlabel metal3 s -960 658052 480 658292 4 io_oeb[24]
port 83 nsew signal tristate
rlabel metal3 s -960 605964 480 606204 4 io_oeb[25]
port 84 nsew signal tristate
rlabel metal3 s -960 553740 480 553980 4 io_oeb[26]
port 85 nsew signal tristate
rlabel metal3 s -960 501652 480 501892 4 io_oeb[27]
port 86 nsew signal tristate
rlabel metal3 s -960 449428 480 449668 4 io_oeb[28]
port 87 nsew signal tristate
rlabel metal3 s -960 397340 480 397580 4 io_oeb[29]
port 88 nsew signal tristate
rlabel metal3 s 583520 112692 584960 112932 6 io_oeb[2]
port 89 nsew signal tristate
rlabel metal3 s -960 345252 480 345492 4 io_oeb[30]
port 90 nsew signal tristate
rlabel metal3 s -960 293028 480 293268 4 io_oeb[31]
port 91 nsew signal tristate
rlabel metal3 s -960 240940 480 241180 4 io_oeb[32]
port 92 nsew signal tristate
rlabel metal3 s -960 188716 480 188956 4 io_oeb[33]
port 93 nsew signal tristate
rlabel metal3 s -960 136628 480 136868 4 io_oeb[34]
port 94 nsew signal tristate
rlabel metal3 s -960 84540 480 84780 4 io_oeb[35]
port 95 nsew signal tristate
rlabel metal3 s -960 45372 480 45612 4 io_oeb[36]
port 96 nsew signal tristate
rlabel metal3 s -960 6340 480 6580 4 io_oeb[37]
port 97 nsew signal tristate
rlabel metal3 s 583520 152540 584960 152780 6 io_oeb[3]
port 98 nsew signal tristate
rlabel metal3 s 583520 192388 584960 192628 6 io_oeb[4]
port 99 nsew signal tristate
rlabel metal3 s 583520 232236 584960 232476 6 io_oeb[5]
port 100 nsew signal tristate
rlabel metal3 s 583520 272084 584960 272324 6 io_oeb[6]
port 101 nsew signal tristate
rlabel metal3 s 583520 325124 584960 325364 6 io_oeb[7]
port 102 nsew signal tristate
rlabel metal3 s 583520 378300 584960 378540 6 io_oeb[8]
port 103 nsew signal tristate
rlabel metal3 s 583520 431476 584960 431716 6 io_oeb[9]
port 104 nsew signal tristate
rlabel metal3 s 583520 19668 584960 19908 6 io_out[0]
port 105 nsew signal tristate
rlabel metal3 s 583520 471324 584960 471564 6 io_out[10]
port 106 nsew signal tristate
rlabel metal3 s 583520 524364 584960 524604 6 io_out[11]
port 107 nsew signal tristate
rlabel metal3 s 583520 577540 584960 577780 6 io_out[12]
port 108 nsew signal tristate
rlabel metal3 s 583520 630716 584960 630956 6 io_out[13]
port 109 nsew signal tristate
rlabel metal3 s 583520 683756 584960 683996 6 io_out[14]
port 110 nsew signal tristate
rlabel metal2 s 543434 703520 543546 704960 6 io_out[15]
port 111 nsew signal tristate
rlabel metal2 s 478482 703520 478594 704960 6 io_out[16]
port 112 nsew signal tristate
rlabel metal2 s 413622 703520 413734 704960 6 io_out[17]
port 113 nsew signal tristate
rlabel metal2 s 348762 703520 348874 704960 6 io_out[18]
port 114 nsew signal tristate
rlabel metal2 s 283810 703520 283922 704960 6 io_out[19]
port 115 nsew signal tristate
rlabel metal3 s 583520 59516 584960 59756 6 io_out[1]
port 116 nsew signal tristate
rlabel metal2 s 218950 703520 219062 704960 6 io_out[20]
port 117 nsew signal tristate
rlabel metal2 s 154090 703520 154202 704960 6 io_out[21]
port 118 nsew signal tristate
rlabel metal2 s 89138 703520 89250 704960 6 io_out[22]
port 119 nsew signal tristate
rlabel metal2 s 24278 703520 24390 704960 6 io_out[23]
port 120 nsew signal tristate
rlabel metal3 s -960 671108 480 671348 4 io_out[24]
port 121 nsew signal tristate
rlabel metal3 s -960 619020 480 619260 4 io_out[25]
port 122 nsew signal tristate
rlabel metal3 s -960 566796 480 567036 4 io_out[26]
port 123 nsew signal tristate
rlabel metal3 s -960 514708 480 514948 4 io_out[27]
port 124 nsew signal tristate
rlabel metal3 s -960 462484 480 462724 4 io_out[28]
port 125 nsew signal tristate
rlabel metal3 s -960 410396 480 410636 4 io_out[29]
port 126 nsew signal tristate
rlabel metal3 s 583520 99364 584960 99604 6 io_out[2]
port 127 nsew signal tristate
rlabel metal3 s -960 358308 480 358548 4 io_out[30]
port 128 nsew signal tristate
rlabel metal3 s -960 306084 480 306324 4 io_out[31]
port 129 nsew signal tristate
rlabel metal3 s -960 253996 480 254236 4 io_out[32]
port 130 nsew signal tristate
rlabel metal3 s -960 201772 480 202012 4 io_out[33]
port 131 nsew signal tristate
rlabel metal3 s -960 149684 480 149924 4 io_out[34]
port 132 nsew signal tristate
rlabel metal3 s -960 97460 480 97700 4 io_out[35]
port 133 nsew signal tristate
rlabel metal3 s -960 58428 480 58668 4 io_out[36]
port 134 nsew signal tristate
rlabel metal3 s -960 19260 480 19500 4 io_out[37]
port 135 nsew signal tristate
rlabel metal3 s 583520 139212 584960 139452 6 io_out[3]
port 136 nsew signal tristate
rlabel metal3 s 583520 179060 584960 179300 6 io_out[4]
port 137 nsew signal tristate
rlabel metal3 s 583520 218908 584960 219148 6 io_out[5]
port 138 nsew signal tristate
rlabel metal3 s 583520 258756 584960 258996 6 io_out[6]
port 139 nsew signal tristate
rlabel metal3 s 583520 311932 584960 312172 6 io_out[7]
port 140 nsew signal tristate
rlabel metal3 s 583520 364972 584960 365212 6 io_out[8]
port 141 nsew signal tristate
rlabel metal3 s 583520 418148 584960 418388 6 io_out[9]
port 142 nsew signal tristate
rlabel metal2 s 125846 -960 125958 480 8 la_data_in[0]
port 143 nsew signal input
rlabel metal2 s 480506 -960 480618 480 8 la_data_in[100]
port 144 nsew signal input
rlabel metal2 s 484002 -960 484114 480 8 la_data_in[101]
port 145 nsew signal input
rlabel metal2 s 487590 -960 487702 480 8 la_data_in[102]
port 146 nsew signal input
rlabel metal2 s 491086 -960 491198 480 8 la_data_in[103]
port 147 nsew signal input
rlabel metal2 s 494674 -960 494786 480 8 la_data_in[104]
port 148 nsew signal input
rlabel metal2 s 498170 -960 498282 480 8 la_data_in[105]
port 149 nsew signal input
rlabel metal2 s 501758 -960 501870 480 8 la_data_in[106]
port 150 nsew signal input
rlabel metal2 s 505346 -960 505458 480 8 la_data_in[107]
port 151 nsew signal input
rlabel metal2 s 508842 -960 508954 480 8 la_data_in[108]
port 152 nsew signal input
rlabel metal2 s 512430 -960 512542 480 8 la_data_in[109]
port 153 nsew signal input
rlabel metal2 s 161266 -960 161378 480 8 la_data_in[10]
port 154 nsew signal input
rlabel metal2 s 515926 -960 516038 480 8 la_data_in[110]
port 155 nsew signal input
rlabel metal2 s 519514 -960 519626 480 8 la_data_in[111]
port 156 nsew signal input
rlabel metal2 s 523010 -960 523122 480 8 la_data_in[112]
port 157 nsew signal input
rlabel metal2 s 526598 -960 526710 480 8 la_data_in[113]
port 158 nsew signal input
rlabel metal2 s 530094 -960 530206 480 8 la_data_in[114]
port 159 nsew signal input
rlabel metal2 s 533682 -960 533794 480 8 la_data_in[115]
port 160 nsew signal input
rlabel metal2 s 537178 -960 537290 480 8 la_data_in[116]
port 161 nsew signal input
rlabel metal2 s 540766 -960 540878 480 8 la_data_in[117]
port 162 nsew signal input
rlabel metal2 s 544354 -960 544466 480 8 la_data_in[118]
port 163 nsew signal input
rlabel metal2 s 547850 -960 547962 480 8 la_data_in[119]
port 164 nsew signal input
rlabel metal2 s 164854 -960 164966 480 8 la_data_in[11]
port 165 nsew signal input
rlabel metal2 s 551438 -960 551550 480 8 la_data_in[120]
port 166 nsew signal input
rlabel metal2 s 554934 -960 555046 480 8 la_data_in[121]
port 167 nsew signal input
rlabel metal2 s 558522 -960 558634 480 8 la_data_in[122]
port 168 nsew signal input
rlabel metal2 s 562018 -960 562130 480 8 la_data_in[123]
port 169 nsew signal input
rlabel metal2 s 565606 -960 565718 480 8 la_data_in[124]
port 170 nsew signal input
rlabel metal2 s 569102 -960 569214 480 8 la_data_in[125]
port 171 nsew signal input
rlabel metal2 s 572690 -960 572802 480 8 la_data_in[126]
port 172 nsew signal input
rlabel metal2 s 576278 -960 576390 480 8 la_data_in[127]
port 173 nsew signal input
rlabel metal2 s 168350 -960 168462 480 8 la_data_in[12]
port 174 nsew signal input
rlabel metal2 s 171938 -960 172050 480 8 la_data_in[13]
port 175 nsew signal input
rlabel metal2 s 175434 -960 175546 480 8 la_data_in[14]
port 176 nsew signal input
rlabel metal2 s 179022 -960 179134 480 8 la_data_in[15]
port 177 nsew signal input
rlabel metal2 s 182518 -960 182630 480 8 la_data_in[16]
port 178 nsew signal input
rlabel metal2 s 186106 -960 186218 480 8 la_data_in[17]
port 179 nsew signal input
rlabel metal2 s 189694 -960 189806 480 8 la_data_in[18]
port 180 nsew signal input
rlabel metal2 s 193190 -960 193302 480 8 la_data_in[19]
port 181 nsew signal input
rlabel metal2 s 129342 -960 129454 480 8 la_data_in[1]
port 182 nsew signal input
rlabel metal2 s 196778 -960 196890 480 8 la_data_in[20]
port 183 nsew signal input
rlabel metal2 s 200274 -960 200386 480 8 la_data_in[21]
port 184 nsew signal input
rlabel metal2 s 203862 -960 203974 480 8 la_data_in[22]
port 185 nsew signal input
rlabel metal2 s 207358 -960 207470 480 8 la_data_in[23]
port 186 nsew signal input
rlabel metal2 s 210946 -960 211058 480 8 la_data_in[24]
port 187 nsew signal input
rlabel metal2 s 214442 -960 214554 480 8 la_data_in[25]
port 188 nsew signal input
rlabel metal2 s 218030 -960 218142 480 8 la_data_in[26]
port 189 nsew signal input
rlabel metal2 s 221526 -960 221638 480 8 la_data_in[27]
port 190 nsew signal input
rlabel metal2 s 225114 -960 225226 480 8 la_data_in[28]
port 191 nsew signal input
rlabel metal2 s 228702 -960 228814 480 8 la_data_in[29]
port 192 nsew signal input
rlabel metal2 s 132930 -960 133042 480 8 la_data_in[2]
port 193 nsew signal input
rlabel metal2 s 232198 -960 232310 480 8 la_data_in[30]
port 194 nsew signal input
rlabel metal2 s 235786 -960 235898 480 8 la_data_in[31]
port 195 nsew signal input
rlabel metal2 s 239282 -960 239394 480 8 la_data_in[32]
port 196 nsew signal input
rlabel metal2 s 242870 -960 242982 480 8 la_data_in[33]
port 197 nsew signal input
rlabel metal2 s 246366 -960 246478 480 8 la_data_in[34]
port 198 nsew signal input
rlabel metal2 s 249954 -960 250066 480 8 la_data_in[35]
port 199 nsew signal input
rlabel metal2 s 253450 -960 253562 480 8 la_data_in[36]
port 200 nsew signal input
rlabel metal2 s 257038 -960 257150 480 8 la_data_in[37]
port 201 nsew signal input
rlabel metal2 s 260626 -960 260738 480 8 la_data_in[38]
port 202 nsew signal input
rlabel metal2 s 264122 -960 264234 480 8 la_data_in[39]
port 203 nsew signal input
rlabel metal2 s 136426 -960 136538 480 8 la_data_in[3]
port 204 nsew signal input
rlabel metal2 s 267710 -960 267822 480 8 la_data_in[40]
port 205 nsew signal input
rlabel metal2 s 271206 -960 271318 480 8 la_data_in[41]
port 206 nsew signal input
rlabel metal2 s 274794 -960 274906 480 8 la_data_in[42]
port 207 nsew signal input
rlabel metal2 s 278290 -960 278402 480 8 la_data_in[43]
port 208 nsew signal input
rlabel metal2 s 281878 -960 281990 480 8 la_data_in[44]
port 209 nsew signal input
rlabel metal2 s 285374 -960 285486 480 8 la_data_in[45]
port 210 nsew signal input
rlabel metal2 s 288962 -960 289074 480 8 la_data_in[46]
port 211 nsew signal input
rlabel metal2 s 292550 -960 292662 480 8 la_data_in[47]
port 212 nsew signal input
rlabel metal2 s 296046 -960 296158 480 8 la_data_in[48]
port 213 nsew signal input
rlabel metal2 s 299634 -960 299746 480 8 la_data_in[49]
port 214 nsew signal input
rlabel metal2 s 140014 -960 140126 480 8 la_data_in[4]
port 215 nsew signal input
rlabel metal2 s 303130 -960 303242 480 8 la_data_in[50]
port 216 nsew signal input
rlabel metal2 s 306718 -960 306830 480 8 la_data_in[51]
port 217 nsew signal input
rlabel metal2 s 310214 -960 310326 480 8 la_data_in[52]
port 218 nsew signal input
rlabel metal2 s 313802 -960 313914 480 8 la_data_in[53]
port 219 nsew signal input
rlabel metal2 s 317298 -960 317410 480 8 la_data_in[54]
port 220 nsew signal input
rlabel metal2 s 320886 -960 320998 480 8 la_data_in[55]
port 221 nsew signal input
rlabel metal2 s 324382 -960 324494 480 8 la_data_in[56]
port 222 nsew signal input
rlabel metal2 s 327970 -960 328082 480 8 la_data_in[57]
port 223 nsew signal input
rlabel metal2 s 331558 -960 331670 480 8 la_data_in[58]
port 224 nsew signal input
rlabel metal2 s 335054 -960 335166 480 8 la_data_in[59]
port 225 nsew signal input
rlabel metal2 s 143510 -960 143622 480 8 la_data_in[5]
port 226 nsew signal input
rlabel metal2 s 338642 -960 338754 480 8 la_data_in[60]
port 227 nsew signal input
rlabel metal2 s 342138 -960 342250 480 8 la_data_in[61]
port 228 nsew signal input
rlabel metal2 s 345726 -960 345838 480 8 la_data_in[62]
port 229 nsew signal input
rlabel metal2 s 349222 -960 349334 480 8 la_data_in[63]
port 230 nsew signal input
rlabel metal2 s 352810 -960 352922 480 8 la_data_in[64]
port 231 nsew signal input
rlabel metal2 s 356306 -960 356418 480 8 la_data_in[65]
port 232 nsew signal input
rlabel metal2 s 359894 -960 360006 480 8 la_data_in[66]
port 233 nsew signal input
rlabel metal2 s 363482 -960 363594 480 8 la_data_in[67]
port 234 nsew signal input
rlabel metal2 s 366978 -960 367090 480 8 la_data_in[68]
port 235 nsew signal input
rlabel metal2 s 370566 -960 370678 480 8 la_data_in[69]
port 236 nsew signal input
rlabel metal2 s 147098 -960 147210 480 8 la_data_in[6]
port 237 nsew signal input
rlabel metal2 s 374062 -960 374174 480 8 la_data_in[70]
port 238 nsew signal input
rlabel metal2 s 377650 -960 377762 480 8 la_data_in[71]
port 239 nsew signal input
rlabel metal2 s 381146 -960 381258 480 8 la_data_in[72]
port 240 nsew signal input
rlabel metal2 s 384734 -960 384846 480 8 la_data_in[73]
port 241 nsew signal input
rlabel metal2 s 388230 -960 388342 480 8 la_data_in[74]
port 242 nsew signal input
rlabel metal2 s 391818 -960 391930 480 8 la_data_in[75]
port 243 nsew signal input
rlabel metal2 s 395314 -960 395426 480 8 la_data_in[76]
port 244 nsew signal input
rlabel metal2 s 398902 -960 399014 480 8 la_data_in[77]
port 245 nsew signal input
rlabel metal2 s 402490 -960 402602 480 8 la_data_in[78]
port 246 nsew signal input
rlabel metal2 s 405986 -960 406098 480 8 la_data_in[79]
port 247 nsew signal input
rlabel metal2 s 150594 -960 150706 480 8 la_data_in[7]
port 248 nsew signal input
rlabel metal2 s 409574 -960 409686 480 8 la_data_in[80]
port 249 nsew signal input
rlabel metal2 s 413070 -960 413182 480 8 la_data_in[81]
port 250 nsew signal input
rlabel metal2 s 416658 -960 416770 480 8 la_data_in[82]
port 251 nsew signal input
rlabel metal2 s 420154 -960 420266 480 8 la_data_in[83]
port 252 nsew signal input
rlabel metal2 s 423742 -960 423854 480 8 la_data_in[84]
port 253 nsew signal input
rlabel metal2 s 427238 -960 427350 480 8 la_data_in[85]
port 254 nsew signal input
rlabel metal2 s 430826 -960 430938 480 8 la_data_in[86]
port 255 nsew signal input
rlabel metal2 s 434414 -960 434526 480 8 la_data_in[87]
port 256 nsew signal input
rlabel metal2 s 437910 -960 438022 480 8 la_data_in[88]
port 257 nsew signal input
rlabel metal2 s 441498 -960 441610 480 8 la_data_in[89]
port 258 nsew signal input
rlabel metal2 s 154182 -960 154294 480 8 la_data_in[8]
port 259 nsew signal input
rlabel metal2 s 444994 -960 445106 480 8 la_data_in[90]
port 260 nsew signal input
rlabel metal2 s 448582 -960 448694 480 8 la_data_in[91]
port 261 nsew signal input
rlabel metal2 s 452078 -960 452190 480 8 la_data_in[92]
port 262 nsew signal input
rlabel metal2 s 455666 -960 455778 480 8 la_data_in[93]
port 263 nsew signal input
rlabel metal2 s 459162 -960 459274 480 8 la_data_in[94]
port 264 nsew signal input
rlabel metal2 s 462750 -960 462862 480 8 la_data_in[95]
port 265 nsew signal input
rlabel metal2 s 466246 -960 466358 480 8 la_data_in[96]
port 266 nsew signal input
rlabel metal2 s 469834 -960 469946 480 8 la_data_in[97]
port 267 nsew signal input
rlabel metal2 s 473422 -960 473534 480 8 la_data_in[98]
port 268 nsew signal input
rlabel metal2 s 476918 -960 477030 480 8 la_data_in[99]
port 269 nsew signal input
rlabel metal2 s 157770 -960 157882 480 8 la_data_in[9]
port 270 nsew signal input
rlabel metal2 s 126950 -960 127062 480 8 la_data_out[0]
port 271 nsew signal tristate
rlabel metal2 s 481702 -960 481814 480 8 la_data_out[100]
port 272 nsew signal tristate
rlabel metal2 s 485198 -960 485310 480 8 la_data_out[101]
port 273 nsew signal tristate
rlabel metal2 s 488786 -960 488898 480 8 la_data_out[102]
port 274 nsew signal tristate
rlabel metal2 s 492282 -960 492394 480 8 la_data_out[103]
port 275 nsew signal tristate
rlabel metal2 s 495870 -960 495982 480 8 la_data_out[104]
port 276 nsew signal tristate
rlabel metal2 s 499366 -960 499478 480 8 la_data_out[105]
port 277 nsew signal tristate
rlabel metal2 s 502954 -960 503066 480 8 la_data_out[106]
port 278 nsew signal tristate
rlabel metal2 s 506450 -960 506562 480 8 la_data_out[107]
port 279 nsew signal tristate
rlabel metal2 s 510038 -960 510150 480 8 la_data_out[108]
port 280 nsew signal tristate
rlabel metal2 s 513534 -960 513646 480 8 la_data_out[109]
port 281 nsew signal tristate
rlabel metal2 s 162462 -960 162574 480 8 la_data_out[10]
port 282 nsew signal tristate
rlabel metal2 s 517122 -960 517234 480 8 la_data_out[110]
port 283 nsew signal tristate
rlabel metal2 s 520710 -960 520822 480 8 la_data_out[111]
port 284 nsew signal tristate
rlabel metal2 s 524206 -960 524318 480 8 la_data_out[112]
port 285 nsew signal tristate
rlabel metal2 s 527794 -960 527906 480 8 la_data_out[113]
port 286 nsew signal tristate
rlabel metal2 s 531290 -960 531402 480 8 la_data_out[114]
port 287 nsew signal tristate
rlabel metal2 s 534878 -960 534990 480 8 la_data_out[115]
port 288 nsew signal tristate
rlabel metal2 s 538374 -960 538486 480 8 la_data_out[116]
port 289 nsew signal tristate
rlabel metal2 s 541962 -960 542074 480 8 la_data_out[117]
port 290 nsew signal tristate
rlabel metal2 s 545458 -960 545570 480 8 la_data_out[118]
port 291 nsew signal tristate
rlabel metal2 s 549046 -960 549158 480 8 la_data_out[119]
port 292 nsew signal tristate
rlabel metal2 s 166050 -960 166162 480 8 la_data_out[11]
port 293 nsew signal tristate
rlabel metal2 s 552634 -960 552746 480 8 la_data_out[120]
port 294 nsew signal tristate
rlabel metal2 s 556130 -960 556242 480 8 la_data_out[121]
port 295 nsew signal tristate
rlabel metal2 s 559718 -960 559830 480 8 la_data_out[122]
port 296 nsew signal tristate
rlabel metal2 s 563214 -960 563326 480 8 la_data_out[123]
port 297 nsew signal tristate
rlabel metal2 s 566802 -960 566914 480 8 la_data_out[124]
port 298 nsew signal tristate
rlabel metal2 s 570298 -960 570410 480 8 la_data_out[125]
port 299 nsew signal tristate
rlabel metal2 s 573886 -960 573998 480 8 la_data_out[126]
port 300 nsew signal tristate
rlabel metal2 s 577382 -960 577494 480 8 la_data_out[127]
port 301 nsew signal tristate
rlabel metal2 s 169546 -960 169658 480 8 la_data_out[12]
port 302 nsew signal tristate
rlabel metal2 s 173134 -960 173246 480 8 la_data_out[13]
port 303 nsew signal tristate
rlabel metal2 s 176630 -960 176742 480 8 la_data_out[14]
port 304 nsew signal tristate
rlabel metal2 s 180218 -960 180330 480 8 la_data_out[15]
port 305 nsew signal tristate
rlabel metal2 s 183714 -960 183826 480 8 la_data_out[16]
port 306 nsew signal tristate
rlabel metal2 s 187302 -960 187414 480 8 la_data_out[17]
port 307 nsew signal tristate
rlabel metal2 s 190798 -960 190910 480 8 la_data_out[18]
port 308 nsew signal tristate
rlabel metal2 s 194386 -960 194498 480 8 la_data_out[19]
port 309 nsew signal tristate
rlabel metal2 s 130538 -960 130650 480 8 la_data_out[1]
port 310 nsew signal tristate
rlabel metal2 s 197882 -960 197994 480 8 la_data_out[20]
port 311 nsew signal tristate
rlabel metal2 s 201470 -960 201582 480 8 la_data_out[21]
port 312 nsew signal tristate
rlabel metal2 s 205058 -960 205170 480 8 la_data_out[22]
port 313 nsew signal tristate
rlabel metal2 s 208554 -960 208666 480 8 la_data_out[23]
port 314 nsew signal tristate
rlabel metal2 s 212142 -960 212254 480 8 la_data_out[24]
port 315 nsew signal tristate
rlabel metal2 s 215638 -960 215750 480 8 la_data_out[25]
port 316 nsew signal tristate
rlabel metal2 s 219226 -960 219338 480 8 la_data_out[26]
port 317 nsew signal tristate
rlabel metal2 s 222722 -960 222834 480 8 la_data_out[27]
port 318 nsew signal tristate
rlabel metal2 s 226310 -960 226422 480 8 la_data_out[28]
port 319 nsew signal tristate
rlabel metal2 s 229806 -960 229918 480 8 la_data_out[29]
port 320 nsew signal tristate
rlabel metal2 s 134126 -960 134238 480 8 la_data_out[2]
port 321 nsew signal tristate
rlabel metal2 s 233394 -960 233506 480 8 la_data_out[30]
port 322 nsew signal tristate
rlabel metal2 s 236982 -960 237094 480 8 la_data_out[31]
port 323 nsew signal tristate
rlabel metal2 s 240478 -960 240590 480 8 la_data_out[32]
port 324 nsew signal tristate
rlabel metal2 s 244066 -960 244178 480 8 la_data_out[33]
port 325 nsew signal tristate
rlabel metal2 s 247562 -960 247674 480 8 la_data_out[34]
port 326 nsew signal tristate
rlabel metal2 s 251150 -960 251262 480 8 la_data_out[35]
port 327 nsew signal tristate
rlabel metal2 s 254646 -960 254758 480 8 la_data_out[36]
port 328 nsew signal tristate
rlabel metal2 s 258234 -960 258346 480 8 la_data_out[37]
port 329 nsew signal tristate
rlabel metal2 s 261730 -960 261842 480 8 la_data_out[38]
port 330 nsew signal tristate
rlabel metal2 s 265318 -960 265430 480 8 la_data_out[39]
port 331 nsew signal tristate
rlabel metal2 s 137622 -960 137734 480 8 la_data_out[3]
port 332 nsew signal tristate
rlabel metal2 s 268814 -960 268926 480 8 la_data_out[40]
port 333 nsew signal tristate
rlabel metal2 s 272402 -960 272514 480 8 la_data_out[41]
port 334 nsew signal tristate
rlabel metal2 s 275990 -960 276102 480 8 la_data_out[42]
port 335 nsew signal tristate
rlabel metal2 s 279486 -960 279598 480 8 la_data_out[43]
port 336 nsew signal tristate
rlabel metal2 s 283074 -960 283186 480 8 la_data_out[44]
port 337 nsew signal tristate
rlabel metal2 s 286570 -960 286682 480 8 la_data_out[45]
port 338 nsew signal tristate
rlabel metal2 s 290158 -960 290270 480 8 la_data_out[46]
port 339 nsew signal tristate
rlabel metal2 s 293654 -960 293766 480 8 la_data_out[47]
port 340 nsew signal tristate
rlabel metal2 s 297242 -960 297354 480 8 la_data_out[48]
port 341 nsew signal tristate
rlabel metal2 s 300738 -960 300850 480 8 la_data_out[49]
port 342 nsew signal tristate
rlabel metal2 s 141210 -960 141322 480 8 la_data_out[4]
port 343 nsew signal tristate
rlabel metal2 s 304326 -960 304438 480 8 la_data_out[50]
port 344 nsew signal tristate
rlabel metal2 s 307914 -960 308026 480 8 la_data_out[51]
port 345 nsew signal tristate
rlabel metal2 s 311410 -960 311522 480 8 la_data_out[52]
port 346 nsew signal tristate
rlabel metal2 s 314998 -960 315110 480 8 la_data_out[53]
port 347 nsew signal tristate
rlabel metal2 s 318494 -960 318606 480 8 la_data_out[54]
port 348 nsew signal tristate
rlabel metal2 s 322082 -960 322194 480 8 la_data_out[55]
port 349 nsew signal tristate
rlabel metal2 s 325578 -960 325690 480 8 la_data_out[56]
port 350 nsew signal tristate
rlabel metal2 s 329166 -960 329278 480 8 la_data_out[57]
port 351 nsew signal tristate
rlabel metal2 s 332662 -960 332774 480 8 la_data_out[58]
port 352 nsew signal tristate
rlabel metal2 s 336250 -960 336362 480 8 la_data_out[59]
port 353 nsew signal tristate
rlabel metal2 s 144706 -960 144818 480 8 la_data_out[5]
port 354 nsew signal tristate
rlabel metal2 s 339838 -960 339950 480 8 la_data_out[60]
port 355 nsew signal tristate
rlabel metal2 s 343334 -960 343446 480 8 la_data_out[61]
port 356 nsew signal tristate
rlabel metal2 s 346922 -960 347034 480 8 la_data_out[62]
port 357 nsew signal tristate
rlabel metal2 s 350418 -960 350530 480 8 la_data_out[63]
port 358 nsew signal tristate
rlabel metal2 s 354006 -960 354118 480 8 la_data_out[64]
port 359 nsew signal tristate
rlabel metal2 s 357502 -960 357614 480 8 la_data_out[65]
port 360 nsew signal tristate
rlabel metal2 s 361090 -960 361202 480 8 la_data_out[66]
port 361 nsew signal tristate
rlabel metal2 s 364586 -960 364698 480 8 la_data_out[67]
port 362 nsew signal tristate
rlabel metal2 s 368174 -960 368286 480 8 la_data_out[68]
port 363 nsew signal tristate
rlabel metal2 s 371670 -960 371782 480 8 la_data_out[69]
port 364 nsew signal tristate
rlabel metal2 s 148294 -960 148406 480 8 la_data_out[6]
port 365 nsew signal tristate
rlabel metal2 s 375258 -960 375370 480 8 la_data_out[70]
port 366 nsew signal tristate
rlabel metal2 s 378846 -960 378958 480 8 la_data_out[71]
port 367 nsew signal tristate
rlabel metal2 s 382342 -960 382454 480 8 la_data_out[72]
port 368 nsew signal tristate
rlabel metal2 s 385930 -960 386042 480 8 la_data_out[73]
port 369 nsew signal tristate
rlabel metal2 s 389426 -960 389538 480 8 la_data_out[74]
port 370 nsew signal tristate
rlabel metal2 s 393014 -960 393126 480 8 la_data_out[75]
port 371 nsew signal tristate
rlabel metal2 s 396510 -960 396622 480 8 la_data_out[76]
port 372 nsew signal tristate
rlabel metal2 s 400098 -960 400210 480 8 la_data_out[77]
port 373 nsew signal tristate
rlabel metal2 s 403594 -960 403706 480 8 la_data_out[78]
port 374 nsew signal tristate
rlabel metal2 s 407182 -960 407294 480 8 la_data_out[79]
port 375 nsew signal tristate
rlabel metal2 s 151790 -960 151902 480 8 la_data_out[7]
port 376 nsew signal tristate
rlabel metal2 s 410770 -960 410882 480 8 la_data_out[80]
port 377 nsew signal tristate
rlabel metal2 s 414266 -960 414378 480 8 la_data_out[81]
port 378 nsew signal tristate
rlabel metal2 s 417854 -960 417966 480 8 la_data_out[82]
port 379 nsew signal tristate
rlabel metal2 s 421350 -960 421462 480 8 la_data_out[83]
port 380 nsew signal tristate
rlabel metal2 s 424938 -960 425050 480 8 la_data_out[84]
port 381 nsew signal tristate
rlabel metal2 s 428434 -960 428546 480 8 la_data_out[85]
port 382 nsew signal tristate
rlabel metal2 s 432022 -960 432134 480 8 la_data_out[86]
port 383 nsew signal tristate
rlabel metal2 s 435518 -960 435630 480 8 la_data_out[87]
port 384 nsew signal tristate
rlabel metal2 s 439106 -960 439218 480 8 la_data_out[88]
port 385 nsew signal tristate
rlabel metal2 s 442602 -960 442714 480 8 la_data_out[89]
port 386 nsew signal tristate
rlabel metal2 s 155378 -960 155490 480 8 la_data_out[8]
port 387 nsew signal tristate
rlabel metal2 s 446190 -960 446302 480 8 la_data_out[90]
port 388 nsew signal tristate
rlabel metal2 s 449778 -960 449890 480 8 la_data_out[91]
port 389 nsew signal tristate
rlabel metal2 s 453274 -960 453386 480 8 la_data_out[92]
port 390 nsew signal tristate
rlabel metal2 s 456862 -960 456974 480 8 la_data_out[93]
port 391 nsew signal tristate
rlabel metal2 s 460358 -960 460470 480 8 la_data_out[94]
port 392 nsew signal tristate
rlabel metal2 s 463946 -960 464058 480 8 la_data_out[95]
port 393 nsew signal tristate
rlabel metal2 s 467442 -960 467554 480 8 la_data_out[96]
port 394 nsew signal tristate
rlabel metal2 s 471030 -960 471142 480 8 la_data_out[97]
port 395 nsew signal tristate
rlabel metal2 s 474526 -960 474638 480 8 la_data_out[98]
port 396 nsew signal tristate
rlabel metal2 s 478114 -960 478226 480 8 la_data_out[99]
port 397 nsew signal tristate
rlabel metal2 s 158874 -960 158986 480 8 la_data_out[9]
port 398 nsew signal tristate
rlabel metal2 s 128146 -960 128258 480 8 la_oenb[0]
port 399 nsew signal input
rlabel metal2 s 482806 -960 482918 480 8 la_oenb[100]
port 400 nsew signal input
rlabel metal2 s 486394 -960 486506 480 8 la_oenb[101]
port 401 nsew signal input
rlabel metal2 s 489890 -960 490002 480 8 la_oenb[102]
port 402 nsew signal input
rlabel metal2 s 493478 -960 493590 480 8 la_oenb[103]
port 403 nsew signal input
rlabel metal2 s 497066 -960 497178 480 8 la_oenb[104]
port 404 nsew signal input
rlabel metal2 s 500562 -960 500674 480 8 la_oenb[105]
port 405 nsew signal input
rlabel metal2 s 504150 -960 504262 480 8 la_oenb[106]
port 406 nsew signal input
rlabel metal2 s 507646 -960 507758 480 8 la_oenb[107]
port 407 nsew signal input
rlabel metal2 s 511234 -960 511346 480 8 la_oenb[108]
port 408 nsew signal input
rlabel metal2 s 514730 -960 514842 480 8 la_oenb[109]
port 409 nsew signal input
rlabel metal2 s 163658 -960 163770 480 8 la_oenb[10]
port 410 nsew signal input
rlabel metal2 s 518318 -960 518430 480 8 la_oenb[110]
port 411 nsew signal input
rlabel metal2 s 521814 -960 521926 480 8 la_oenb[111]
port 412 nsew signal input
rlabel metal2 s 525402 -960 525514 480 8 la_oenb[112]
port 413 nsew signal input
rlabel metal2 s 528990 -960 529102 480 8 la_oenb[113]
port 414 nsew signal input
rlabel metal2 s 532486 -960 532598 480 8 la_oenb[114]
port 415 nsew signal input
rlabel metal2 s 536074 -960 536186 480 8 la_oenb[115]
port 416 nsew signal input
rlabel metal2 s 539570 -960 539682 480 8 la_oenb[116]
port 417 nsew signal input
rlabel metal2 s 543158 -960 543270 480 8 la_oenb[117]
port 418 nsew signal input
rlabel metal2 s 546654 -960 546766 480 8 la_oenb[118]
port 419 nsew signal input
rlabel metal2 s 550242 -960 550354 480 8 la_oenb[119]
port 420 nsew signal input
rlabel metal2 s 167154 -960 167266 480 8 la_oenb[11]
port 421 nsew signal input
rlabel metal2 s 553738 -960 553850 480 8 la_oenb[120]
port 422 nsew signal input
rlabel metal2 s 557326 -960 557438 480 8 la_oenb[121]
port 423 nsew signal input
rlabel metal2 s 560822 -960 560934 480 8 la_oenb[122]
port 424 nsew signal input
rlabel metal2 s 564410 -960 564522 480 8 la_oenb[123]
port 425 nsew signal input
rlabel metal2 s 567998 -960 568110 480 8 la_oenb[124]
port 426 nsew signal input
rlabel metal2 s 571494 -960 571606 480 8 la_oenb[125]
port 427 nsew signal input
rlabel metal2 s 575082 -960 575194 480 8 la_oenb[126]
port 428 nsew signal input
rlabel metal2 s 578578 -960 578690 480 8 la_oenb[127]
port 429 nsew signal input
rlabel metal2 s 170742 -960 170854 480 8 la_oenb[12]
port 430 nsew signal input
rlabel metal2 s 174238 -960 174350 480 8 la_oenb[13]
port 431 nsew signal input
rlabel metal2 s 177826 -960 177938 480 8 la_oenb[14]
port 432 nsew signal input
rlabel metal2 s 181414 -960 181526 480 8 la_oenb[15]
port 433 nsew signal input
rlabel metal2 s 184910 -960 185022 480 8 la_oenb[16]
port 434 nsew signal input
rlabel metal2 s 188498 -960 188610 480 8 la_oenb[17]
port 435 nsew signal input
rlabel metal2 s 191994 -960 192106 480 8 la_oenb[18]
port 436 nsew signal input
rlabel metal2 s 195582 -960 195694 480 8 la_oenb[19]
port 437 nsew signal input
rlabel metal2 s 131734 -960 131846 480 8 la_oenb[1]
port 438 nsew signal input
rlabel metal2 s 199078 -960 199190 480 8 la_oenb[20]
port 439 nsew signal input
rlabel metal2 s 202666 -960 202778 480 8 la_oenb[21]
port 440 nsew signal input
rlabel metal2 s 206162 -960 206274 480 8 la_oenb[22]
port 441 nsew signal input
rlabel metal2 s 209750 -960 209862 480 8 la_oenb[23]
port 442 nsew signal input
rlabel metal2 s 213338 -960 213450 480 8 la_oenb[24]
port 443 nsew signal input
rlabel metal2 s 216834 -960 216946 480 8 la_oenb[25]
port 444 nsew signal input
rlabel metal2 s 220422 -960 220534 480 8 la_oenb[26]
port 445 nsew signal input
rlabel metal2 s 223918 -960 224030 480 8 la_oenb[27]
port 446 nsew signal input
rlabel metal2 s 227506 -960 227618 480 8 la_oenb[28]
port 447 nsew signal input
rlabel metal2 s 231002 -960 231114 480 8 la_oenb[29]
port 448 nsew signal input
rlabel metal2 s 135230 -960 135342 480 8 la_oenb[2]
port 449 nsew signal input
rlabel metal2 s 234590 -960 234702 480 8 la_oenb[30]
port 450 nsew signal input
rlabel metal2 s 238086 -960 238198 480 8 la_oenb[31]
port 451 nsew signal input
rlabel metal2 s 241674 -960 241786 480 8 la_oenb[32]
port 452 nsew signal input
rlabel metal2 s 245170 -960 245282 480 8 la_oenb[33]
port 453 nsew signal input
rlabel metal2 s 248758 -960 248870 480 8 la_oenb[34]
port 454 nsew signal input
rlabel metal2 s 252346 -960 252458 480 8 la_oenb[35]
port 455 nsew signal input
rlabel metal2 s 255842 -960 255954 480 8 la_oenb[36]
port 456 nsew signal input
rlabel metal2 s 259430 -960 259542 480 8 la_oenb[37]
port 457 nsew signal input
rlabel metal2 s 262926 -960 263038 480 8 la_oenb[38]
port 458 nsew signal input
rlabel metal2 s 266514 -960 266626 480 8 la_oenb[39]
port 459 nsew signal input
rlabel metal2 s 138818 -960 138930 480 8 la_oenb[3]
port 460 nsew signal input
rlabel metal2 s 270010 -960 270122 480 8 la_oenb[40]
port 461 nsew signal input
rlabel metal2 s 273598 -960 273710 480 8 la_oenb[41]
port 462 nsew signal input
rlabel metal2 s 277094 -960 277206 480 8 la_oenb[42]
port 463 nsew signal input
rlabel metal2 s 280682 -960 280794 480 8 la_oenb[43]
port 464 nsew signal input
rlabel metal2 s 284270 -960 284382 480 8 la_oenb[44]
port 465 nsew signal input
rlabel metal2 s 287766 -960 287878 480 8 la_oenb[45]
port 466 nsew signal input
rlabel metal2 s 291354 -960 291466 480 8 la_oenb[46]
port 467 nsew signal input
rlabel metal2 s 294850 -960 294962 480 8 la_oenb[47]
port 468 nsew signal input
rlabel metal2 s 298438 -960 298550 480 8 la_oenb[48]
port 469 nsew signal input
rlabel metal2 s 301934 -960 302046 480 8 la_oenb[49]
port 470 nsew signal input
rlabel metal2 s 142406 -960 142518 480 8 la_oenb[4]
port 471 nsew signal input
rlabel metal2 s 305522 -960 305634 480 8 la_oenb[50]
port 472 nsew signal input
rlabel metal2 s 309018 -960 309130 480 8 la_oenb[51]
port 473 nsew signal input
rlabel metal2 s 312606 -960 312718 480 8 la_oenb[52]
port 474 nsew signal input
rlabel metal2 s 316194 -960 316306 480 8 la_oenb[53]
port 475 nsew signal input
rlabel metal2 s 319690 -960 319802 480 8 la_oenb[54]
port 476 nsew signal input
rlabel metal2 s 323278 -960 323390 480 8 la_oenb[55]
port 477 nsew signal input
rlabel metal2 s 326774 -960 326886 480 8 la_oenb[56]
port 478 nsew signal input
rlabel metal2 s 330362 -960 330474 480 8 la_oenb[57]
port 479 nsew signal input
rlabel metal2 s 333858 -960 333970 480 8 la_oenb[58]
port 480 nsew signal input
rlabel metal2 s 337446 -960 337558 480 8 la_oenb[59]
port 481 nsew signal input
rlabel metal2 s 145902 -960 146014 480 8 la_oenb[5]
port 482 nsew signal input
rlabel metal2 s 340942 -960 341054 480 8 la_oenb[60]
port 483 nsew signal input
rlabel metal2 s 344530 -960 344642 480 8 la_oenb[61]
port 484 nsew signal input
rlabel metal2 s 348026 -960 348138 480 8 la_oenb[62]
port 485 nsew signal input
rlabel metal2 s 351614 -960 351726 480 8 la_oenb[63]
port 486 nsew signal input
rlabel metal2 s 355202 -960 355314 480 8 la_oenb[64]
port 487 nsew signal input
rlabel metal2 s 358698 -960 358810 480 8 la_oenb[65]
port 488 nsew signal input
rlabel metal2 s 362286 -960 362398 480 8 la_oenb[66]
port 489 nsew signal input
rlabel metal2 s 365782 -960 365894 480 8 la_oenb[67]
port 490 nsew signal input
rlabel metal2 s 369370 -960 369482 480 8 la_oenb[68]
port 491 nsew signal input
rlabel metal2 s 372866 -960 372978 480 8 la_oenb[69]
port 492 nsew signal input
rlabel metal2 s 149490 -960 149602 480 8 la_oenb[6]
port 493 nsew signal input
rlabel metal2 s 376454 -960 376566 480 8 la_oenb[70]
port 494 nsew signal input
rlabel metal2 s 379950 -960 380062 480 8 la_oenb[71]
port 495 nsew signal input
rlabel metal2 s 383538 -960 383650 480 8 la_oenb[72]
port 496 nsew signal input
rlabel metal2 s 387126 -960 387238 480 8 la_oenb[73]
port 497 nsew signal input
rlabel metal2 s 390622 -960 390734 480 8 la_oenb[74]
port 498 nsew signal input
rlabel metal2 s 394210 -960 394322 480 8 la_oenb[75]
port 499 nsew signal input
rlabel metal2 s 397706 -960 397818 480 8 la_oenb[76]
port 500 nsew signal input
rlabel metal2 s 401294 -960 401406 480 8 la_oenb[77]
port 501 nsew signal input
rlabel metal2 s 404790 -960 404902 480 8 la_oenb[78]
port 502 nsew signal input
rlabel metal2 s 408378 -960 408490 480 8 la_oenb[79]
port 503 nsew signal input
rlabel metal2 s 152986 -960 153098 480 8 la_oenb[7]
port 504 nsew signal input
rlabel metal2 s 411874 -960 411986 480 8 la_oenb[80]
port 505 nsew signal input
rlabel metal2 s 415462 -960 415574 480 8 la_oenb[81]
port 506 nsew signal input
rlabel metal2 s 418958 -960 419070 480 8 la_oenb[82]
port 507 nsew signal input
rlabel metal2 s 422546 -960 422658 480 8 la_oenb[83]
port 508 nsew signal input
rlabel metal2 s 426134 -960 426246 480 8 la_oenb[84]
port 509 nsew signal input
rlabel metal2 s 429630 -960 429742 480 8 la_oenb[85]
port 510 nsew signal input
rlabel metal2 s 433218 -960 433330 480 8 la_oenb[86]
port 511 nsew signal input
rlabel metal2 s 436714 -960 436826 480 8 la_oenb[87]
port 512 nsew signal input
rlabel metal2 s 440302 -960 440414 480 8 la_oenb[88]
port 513 nsew signal input
rlabel metal2 s 443798 -960 443910 480 8 la_oenb[89]
port 514 nsew signal input
rlabel metal2 s 156574 -960 156686 480 8 la_oenb[8]
port 515 nsew signal input
rlabel metal2 s 447386 -960 447498 480 8 la_oenb[90]
port 516 nsew signal input
rlabel metal2 s 450882 -960 450994 480 8 la_oenb[91]
port 517 nsew signal input
rlabel metal2 s 454470 -960 454582 480 8 la_oenb[92]
port 518 nsew signal input
rlabel metal2 s 458058 -960 458170 480 8 la_oenb[93]
port 519 nsew signal input
rlabel metal2 s 461554 -960 461666 480 8 la_oenb[94]
port 520 nsew signal input
rlabel metal2 s 465142 -960 465254 480 8 la_oenb[95]
port 521 nsew signal input
rlabel metal2 s 468638 -960 468750 480 8 la_oenb[96]
port 522 nsew signal input
rlabel metal2 s 472226 -960 472338 480 8 la_oenb[97]
port 523 nsew signal input
rlabel metal2 s 475722 -960 475834 480 8 la_oenb[98]
port 524 nsew signal input
rlabel metal2 s 479310 -960 479422 480 8 la_oenb[99]
port 525 nsew signal input
rlabel metal2 s 160070 -960 160182 480 8 la_oenb[9]
port 526 nsew signal input
rlabel metal2 s 579774 -960 579886 480 8 user_clock2
port 527 nsew signal input
rlabel metal2 s 580970 -960 581082 480 8 user_irq[0]
port 528 nsew signal tristate
rlabel metal2 s 582166 -960 582278 480 8 user_irq[1]
port 529 nsew signal tristate
rlabel metal2 s 583362 -960 583474 480 8 user_irq[2]
port 530 nsew signal tristate
rlabel metal5 s -2006 -934 585930 -314 8 vccd1
port 531 nsew power input
rlabel metal5 s -2966 1876 586890 2476 6 vccd1
port 531 nsew power input
rlabel metal5 s -2966 37876 586890 38476 6 vccd1
port 531 nsew power input
rlabel metal5 s -2966 73876 586890 74476 6 vccd1
port 531 nsew power input
rlabel metal5 s -2966 109876 586890 110476 6 vccd1
port 531 nsew power input
rlabel metal5 s -2966 145876 586890 146476 6 vccd1
port 531 nsew power input
rlabel metal5 s -2966 181876 586890 182476 6 vccd1
port 531 nsew power input
rlabel metal5 s -2966 217876 586890 218476 6 vccd1
port 531 nsew power input
rlabel metal5 s -2966 253876 586890 254476 6 vccd1
port 531 nsew power input
rlabel metal5 s -2966 289876 586890 290476 6 vccd1
port 531 nsew power input
rlabel metal5 s -2966 325876 586890 326476 6 vccd1
port 531 nsew power input
rlabel metal5 s -2966 361876 586890 362476 6 vccd1
port 531 nsew power input
rlabel metal5 s -2966 397876 586890 398476 6 vccd1
port 531 nsew power input
rlabel metal5 s -2966 433876 586890 434476 6 vccd1
port 531 nsew power input
rlabel metal5 s -2966 469876 586890 470476 6 vccd1
port 531 nsew power input
rlabel metal5 s -2966 505876 586890 506476 6 vccd1
port 531 nsew power input
rlabel metal5 s -2966 541876 586890 542476 6 vccd1
port 531 nsew power input
rlabel metal5 s -2966 577876 586890 578476 6 vccd1
port 531 nsew power input
rlabel metal5 s -2966 613876 586890 614476 6 vccd1
port 531 nsew power input
rlabel metal5 s -2966 649876 586890 650476 6 vccd1
port 531 nsew power input
rlabel metal5 s -2966 685876 586890 686476 6 vccd1
port 531 nsew power input
rlabel metal5 s -2006 704250 585930 704870 6 vccd1
port 531 nsew power input
rlabel metal4 s 72804 -1894 73404 38000 6 vccd1
port 531 nsew power input
rlabel metal4 s 108804 -1894 109404 38000 6 vccd1
port 531 nsew power input
rlabel metal4 s 144804 -1894 145404 38000 6 vccd1
port 531 nsew power input
rlabel metal4 s 180804 -1894 181404 38000 6 vccd1
port 531 nsew power input
rlabel metal4 s 216804 -1894 217404 38000 6 vccd1
port 531 nsew power input
rlabel metal4 s 72804 242304 73404 338000 6 vccd1
port 531 nsew power input
rlabel metal4 s 108804 242304 109404 338000 6 vccd1
port 531 nsew power input
rlabel metal4 s 144804 242304 145404 338000 6 vccd1
port 531 nsew power input
rlabel metal4 s 360804 -1894 361404 338000 6 vccd1
port 531 nsew power input
rlabel metal4 s 396804 -1894 397404 338000 6 vccd1
port 531 nsew power input
rlabel metal4 s 432804 -1894 433404 338000 6 vccd1
port 531 nsew power input
rlabel metal4 s 468804 -1894 469404 338000 6 vccd1
port 531 nsew power input
rlabel metal4 s -2006 -934 -1386 704870 4 vccd1
port 531 nsew power input
rlabel metal4 s 585310 -934 585930 704870 6 vccd1
port 531 nsew power input
rlabel metal4 s 804 -1894 1404 705830 6 vccd1
port 531 nsew power input
rlabel metal4 s 36804 -1894 37404 705830 6 vccd1
port 531 nsew power input
rlabel metal4 s 72804 425308 73404 705830 6 vccd1
port 531 nsew power input
rlabel metal4 s 108804 425308 109404 705830 6 vccd1
port 531 nsew power input
rlabel metal4 s 144804 425308 145404 705830 6 vccd1
port 531 nsew power input
rlabel metal4 s 180804 242304 181404 705830 6 vccd1
port 531 nsew power input
rlabel metal4 s 216804 242304 217404 705830 6 vccd1
port 531 nsew power input
rlabel metal4 s 252804 -1894 253404 705830 6 vccd1
port 531 nsew power input
rlabel metal4 s 288804 -1894 289404 705830 6 vccd1
port 531 nsew power input
rlabel metal4 s 324804 -1894 325404 705830 6 vccd1
port 531 nsew power input
rlabel metal4 s 360804 425308 361404 705830 6 vccd1
port 531 nsew power input
rlabel metal4 s 396804 425308 397404 705830 6 vccd1
port 531 nsew power input
rlabel metal4 s 432804 425308 433404 705830 6 vccd1
port 531 nsew power input
rlabel metal4 s 468804 425308 469404 705830 6 vccd1
port 531 nsew power input
rlabel metal4 s 504804 -1894 505404 705830 6 vccd1
port 531 nsew power input
rlabel metal4 s 540804 -1894 541404 705830 6 vccd1
port 531 nsew power input
rlabel metal4 s 576804 -1894 577404 705830 6 vccd1
port 531 nsew power input
rlabel metal5 s -3926 -2854 587850 -2234 8 vccd2
port 532 nsew power input
rlabel metal5 s -4886 5576 588810 6176 6 vccd2
port 532 nsew power input
rlabel metal5 s -4886 41576 588810 42176 6 vccd2
port 532 nsew power input
rlabel metal5 s -4886 77576 588810 78176 6 vccd2
port 532 nsew power input
rlabel metal5 s -4886 113576 588810 114176 6 vccd2
port 532 nsew power input
rlabel metal5 s -4886 149576 588810 150176 6 vccd2
port 532 nsew power input
rlabel metal5 s -4886 185576 588810 186176 6 vccd2
port 532 nsew power input
rlabel metal5 s -4886 221576 588810 222176 6 vccd2
port 532 nsew power input
rlabel metal5 s -4886 257576 588810 258176 6 vccd2
port 532 nsew power input
rlabel metal5 s -4886 293576 588810 294176 6 vccd2
port 532 nsew power input
rlabel metal5 s -4886 329576 588810 330176 6 vccd2
port 532 nsew power input
rlabel metal5 s -4886 365576 588810 366176 6 vccd2
port 532 nsew power input
rlabel metal5 s -4886 401576 588810 402176 6 vccd2
port 532 nsew power input
rlabel metal5 s -4886 437576 588810 438176 6 vccd2
port 532 nsew power input
rlabel metal5 s -4886 473576 588810 474176 6 vccd2
port 532 nsew power input
rlabel metal5 s -4886 509576 588810 510176 6 vccd2
port 532 nsew power input
rlabel metal5 s -4886 545576 588810 546176 6 vccd2
port 532 nsew power input
rlabel metal5 s -4886 581576 588810 582176 6 vccd2
port 532 nsew power input
rlabel metal5 s -4886 617576 588810 618176 6 vccd2
port 532 nsew power input
rlabel metal5 s -4886 653576 588810 654176 6 vccd2
port 532 nsew power input
rlabel metal5 s -4886 689576 588810 690176 6 vccd2
port 532 nsew power input
rlabel metal5 s -3926 706170 587850 706790 6 vccd2
port 532 nsew power input
rlabel metal4 s 40504 -3814 41104 38000 6 vccd2
port 532 nsew power input
rlabel metal4 s 76504 -3814 77104 38000 6 vccd2
port 532 nsew power input
rlabel metal4 s 112504 -3814 113104 38000 6 vccd2
port 532 nsew power input
rlabel metal4 s 148504 -3814 149104 38000 6 vccd2
port 532 nsew power input
rlabel metal4 s 184504 -3814 185104 38000 6 vccd2
port 532 nsew power input
rlabel metal4 s 220504 -3814 221104 38000 6 vccd2
port 532 nsew power input
rlabel metal4 s 40504 242304 41104 338000 6 vccd2
port 532 nsew power input
rlabel metal4 s 76504 242304 77104 338000 6 vccd2
port 532 nsew power input
rlabel metal4 s 112504 242304 113104 338000 6 vccd2
port 532 nsew power input
rlabel metal4 s 148504 242304 149104 338000 6 vccd2
port 532 nsew power input
rlabel metal4 s 364504 -3814 365104 338000 6 vccd2
port 532 nsew power input
rlabel metal4 s 400504 -3814 401104 338000 6 vccd2
port 532 nsew power input
rlabel metal4 s 436504 -3814 437104 338000 6 vccd2
port 532 nsew power input
rlabel metal4 s 472504 -3814 473104 338000 6 vccd2
port 532 nsew power input
rlabel metal4 s -3926 -2854 -3306 706790 4 vccd2
port 532 nsew power input
rlabel metal4 s 587230 -2854 587850 706790 6 vccd2
port 532 nsew power input
rlabel metal4 s 4504 -3814 5104 707750 6 vccd2
port 532 nsew power input
rlabel metal4 s 40504 425308 41104 707750 6 vccd2
port 532 nsew power input
rlabel metal4 s 76504 425308 77104 707750 6 vccd2
port 532 nsew power input
rlabel metal4 s 112504 425308 113104 707750 6 vccd2
port 532 nsew power input
rlabel metal4 s 148504 425308 149104 707750 6 vccd2
port 532 nsew power input
rlabel metal4 s 184504 242304 185104 707750 6 vccd2
port 532 nsew power input
rlabel metal4 s 220504 242304 221104 707750 6 vccd2
port 532 nsew power input
rlabel metal4 s 256504 -3814 257104 707750 6 vccd2
port 532 nsew power input
rlabel metal4 s 292504 -3814 293104 707750 6 vccd2
port 532 nsew power input
rlabel metal4 s 328504 -3814 329104 707750 6 vccd2
port 532 nsew power input
rlabel metal4 s 364504 425308 365104 707750 6 vccd2
port 532 nsew power input
rlabel metal4 s 400504 425308 401104 707750 6 vccd2
port 532 nsew power input
rlabel metal4 s 436504 425308 437104 707750 6 vccd2
port 532 nsew power input
rlabel metal4 s 472504 425308 473104 707750 6 vccd2
port 532 nsew power input
rlabel metal4 s 508504 -3814 509104 707750 6 vccd2
port 532 nsew power input
rlabel metal4 s 544504 -3814 545104 707750 6 vccd2
port 532 nsew power input
rlabel metal4 s 580504 -3814 581104 707750 6 vccd2
port 532 nsew power input
rlabel metal5 s -5846 -4774 589770 -4154 8 vdda1
port 533 nsew power input
rlabel metal5 s -6806 9276 590730 9876 6 vdda1
port 533 nsew power input
rlabel metal5 s -6806 45276 590730 45876 6 vdda1
port 533 nsew power input
rlabel metal5 s -6806 81276 590730 81876 6 vdda1
port 533 nsew power input
rlabel metal5 s -6806 117276 590730 117876 6 vdda1
port 533 nsew power input
rlabel metal5 s -6806 153276 590730 153876 6 vdda1
port 533 nsew power input
rlabel metal5 s -6806 189276 590730 189876 6 vdda1
port 533 nsew power input
rlabel metal5 s -6806 225276 590730 225876 6 vdda1
port 533 nsew power input
rlabel metal5 s -6806 261276 590730 261876 6 vdda1
port 533 nsew power input
rlabel metal5 s -6806 297276 590730 297876 6 vdda1
port 533 nsew power input
rlabel metal5 s -6806 333276 590730 333876 6 vdda1
port 533 nsew power input
rlabel metal5 s -6806 369276 590730 369876 6 vdda1
port 533 nsew power input
rlabel metal5 s -6806 405276 590730 405876 6 vdda1
port 533 nsew power input
rlabel metal5 s -6806 441276 590730 441876 6 vdda1
port 533 nsew power input
rlabel metal5 s -6806 477276 590730 477876 6 vdda1
port 533 nsew power input
rlabel metal5 s -6806 513276 590730 513876 6 vdda1
port 533 nsew power input
rlabel metal5 s -6806 549276 590730 549876 6 vdda1
port 533 nsew power input
rlabel metal5 s -6806 585276 590730 585876 6 vdda1
port 533 nsew power input
rlabel metal5 s -6806 621276 590730 621876 6 vdda1
port 533 nsew power input
rlabel metal5 s -6806 657276 590730 657876 6 vdda1
port 533 nsew power input
rlabel metal5 s -6806 693276 590730 693876 6 vdda1
port 533 nsew power input
rlabel metal5 s -5846 708090 589770 708710 6 vdda1
port 533 nsew power input
rlabel metal4 s 44204 -5734 44804 38000 6 vdda1
port 533 nsew power input
rlabel metal4 s 80204 -5734 80804 38000 6 vdda1
port 533 nsew power input
rlabel metal4 s 116204 -5734 116804 38000 6 vdda1
port 533 nsew power input
rlabel metal4 s 152204 -5734 152804 38000 6 vdda1
port 533 nsew power input
rlabel metal4 s 188204 -5734 188804 38000 6 vdda1
port 533 nsew power input
rlabel metal4 s 224204 -5734 224804 38000 6 vdda1
port 533 nsew power input
rlabel metal4 s 44204 242304 44804 338000 6 vdda1
port 533 nsew power input
rlabel metal4 s 80204 242304 80804 338000 6 vdda1
port 533 nsew power input
rlabel metal4 s 116204 242304 116804 338000 6 vdda1
port 533 nsew power input
rlabel metal4 s 152204 242304 152804 338000 6 vdda1
port 533 nsew power input
rlabel metal4 s 368204 -5734 368804 338000 6 vdda1
port 533 nsew power input
rlabel metal4 s 404204 -5734 404804 338000 6 vdda1
port 533 nsew power input
rlabel metal4 s 440204 -5734 440804 338000 6 vdda1
port 533 nsew power input
rlabel metal4 s 476204 -5734 476804 338000 6 vdda1
port 533 nsew power input
rlabel metal4 s -5846 -4774 -5226 708710 4 vdda1
port 533 nsew power input
rlabel metal4 s 589150 -4774 589770 708710 6 vdda1
port 533 nsew power input
rlabel metal4 s 8204 -5734 8804 709670 6 vdda1
port 533 nsew power input
rlabel metal4 s 44204 425308 44804 709670 6 vdda1
port 533 nsew power input
rlabel metal4 s 80204 425308 80804 709670 6 vdda1
port 533 nsew power input
rlabel metal4 s 116204 425308 116804 709670 6 vdda1
port 533 nsew power input
rlabel metal4 s 152204 425308 152804 709670 6 vdda1
port 533 nsew power input
rlabel metal4 s 188204 242304 188804 709670 6 vdda1
port 533 nsew power input
rlabel metal4 s 224204 242304 224804 709670 6 vdda1
port 533 nsew power input
rlabel metal4 s 260204 -5734 260804 709670 6 vdda1
port 533 nsew power input
rlabel metal4 s 296204 -5734 296804 709670 6 vdda1
port 533 nsew power input
rlabel metal4 s 332204 -5734 332804 709670 6 vdda1
port 533 nsew power input
rlabel metal4 s 368204 425308 368804 709670 6 vdda1
port 533 nsew power input
rlabel metal4 s 404204 425308 404804 709670 6 vdda1
port 533 nsew power input
rlabel metal4 s 440204 425308 440804 709670 6 vdda1
port 533 nsew power input
rlabel metal4 s 476204 425308 476804 709670 6 vdda1
port 533 nsew power input
rlabel metal4 s 512204 -5734 512804 709670 6 vdda1
port 533 nsew power input
rlabel metal4 s 548204 -5734 548804 709670 6 vdda1
port 533 nsew power input
rlabel metal5 s -7766 -6694 591690 -6074 8 vdda2
port 534 nsew power input
rlabel metal5 s -8726 12976 592650 13576 6 vdda2
port 534 nsew power input
rlabel metal5 s -8726 48976 592650 49576 6 vdda2
port 534 nsew power input
rlabel metal5 s -8726 84976 592650 85576 6 vdda2
port 534 nsew power input
rlabel metal5 s -8726 120976 592650 121576 6 vdda2
port 534 nsew power input
rlabel metal5 s -8726 156976 592650 157576 6 vdda2
port 534 nsew power input
rlabel metal5 s -8726 192976 592650 193576 6 vdda2
port 534 nsew power input
rlabel metal5 s -8726 228976 592650 229576 6 vdda2
port 534 nsew power input
rlabel metal5 s -8726 264976 592650 265576 6 vdda2
port 534 nsew power input
rlabel metal5 s -8726 300976 592650 301576 6 vdda2
port 534 nsew power input
rlabel metal5 s -8726 336976 592650 337576 6 vdda2
port 534 nsew power input
rlabel metal5 s -8726 372976 592650 373576 6 vdda2
port 534 nsew power input
rlabel metal5 s -8726 408976 592650 409576 6 vdda2
port 534 nsew power input
rlabel metal5 s -8726 444976 592650 445576 6 vdda2
port 534 nsew power input
rlabel metal5 s -8726 480976 592650 481576 6 vdda2
port 534 nsew power input
rlabel metal5 s -8726 516976 592650 517576 6 vdda2
port 534 nsew power input
rlabel metal5 s -8726 552976 592650 553576 6 vdda2
port 534 nsew power input
rlabel metal5 s -8726 588976 592650 589576 6 vdda2
port 534 nsew power input
rlabel metal5 s -8726 624976 592650 625576 6 vdda2
port 534 nsew power input
rlabel metal5 s -8726 660976 592650 661576 6 vdda2
port 534 nsew power input
rlabel metal5 s -8726 696976 592650 697576 6 vdda2
port 534 nsew power input
rlabel metal5 s -7766 710010 591690 710630 6 vdda2
port 534 nsew power input
rlabel metal4 s 47904 -7654 48504 38000 6 vdda2
port 534 nsew power input
rlabel metal4 s 83904 -7654 84504 38000 6 vdda2
port 534 nsew power input
rlabel metal4 s 119904 -7654 120504 38000 6 vdda2
port 534 nsew power input
rlabel metal4 s 155904 -7654 156504 38000 6 vdda2
port 534 nsew power input
rlabel metal4 s 191904 -7654 192504 38000 6 vdda2
port 534 nsew power input
rlabel metal4 s 227904 -7654 228504 38000 6 vdda2
port 534 nsew power input
rlabel metal4 s 47904 242304 48504 338000 6 vdda2
port 534 nsew power input
rlabel metal4 s 83904 242304 84504 338000 6 vdda2
port 534 nsew power input
rlabel metal4 s 119904 242304 120504 338000 6 vdda2
port 534 nsew power input
rlabel metal4 s 155904 242304 156504 338000 6 vdda2
port 534 nsew power input
rlabel metal4 s 371904 -7654 372504 338000 6 vdda2
port 534 nsew power input
rlabel metal4 s 407904 -7654 408504 338000 6 vdda2
port 534 nsew power input
rlabel metal4 s 443904 -7654 444504 338000 6 vdda2
port 534 nsew power input
rlabel metal4 s -7766 -6694 -7146 710630 4 vdda2
port 534 nsew power input
rlabel metal4 s 591070 -6694 591690 710630 6 vdda2
port 534 nsew power input
rlabel metal4 s 11904 -7654 12504 711590 6 vdda2
port 534 nsew power input
rlabel metal4 s 47904 425308 48504 711590 6 vdda2
port 534 nsew power input
rlabel metal4 s 83904 425308 84504 711590 6 vdda2
port 534 nsew power input
rlabel metal4 s 119904 425308 120504 711590 6 vdda2
port 534 nsew power input
rlabel metal4 s 155904 425308 156504 711590 6 vdda2
port 534 nsew power input
rlabel metal4 s 191904 242304 192504 711590 6 vdda2
port 534 nsew power input
rlabel metal4 s 227904 242304 228504 711590 6 vdda2
port 534 nsew power input
rlabel metal4 s 263904 -7654 264504 711590 6 vdda2
port 534 nsew power input
rlabel metal4 s 299904 -7654 300504 711590 6 vdda2
port 534 nsew power input
rlabel metal4 s 335904 -7654 336504 711590 6 vdda2
port 534 nsew power input
rlabel metal4 s 371904 425308 372504 711590 6 vdda2
port 534 nsew power input
rlabel metal4 s 407904 425308 408504 711590 6 vdda2
port 534 nsew power input
rlabel metal4 s 443904 425308 444504 711590 6 vdda2
port 534 nsew power input
rlabel metal4 s 479904 -7654 480504 711590 6 vdda2
port 534 nsew power input
rlabel metal4 s 515904 -7654 516504 711590 6 vdda2
port 534 nsew power input
rlabel metal4 s 551904 -7654 552504 711590 6 vdda2
port 534 nsew power input
rlabel metal5 s -6806 -5734 590730 -5114 8 vssa1
port 535 nsew ground input
rlabel metal5 s -6806 27276 590730 27876 6 vssa1
port 535 nsew ground input
rlabel metal5 s -6806 63276 590730 63876 6 vssa1
port 535 nsew ground input
rlabel metal5 s -6806 99276 590730 99876 6 vssa1
port 535 nsew ground input
rlabel metal5 s -6806 135276 590730 135876 6 vssa1
port 535 nsew ground input
rlabel metal5 s -6806 171276 590730 171876 6 vssa1
port 535 nsew ground input
rlabel metal5 s -6806 207276 590730 207876 6 vssa1
port 535 nsew ground input
rlabel metal5 s -6806 243276 590730 243876 6 vssa1
port 535 nsew ground input
rlabel metal5 s -6806 279276 590730 279876 6 vssa1
port 535 nsew ground input
rlabel metal5 s -6806 315276 590730 315876 6 vssa1
port 535 nsew ground input
rlabel metal5 s -6806 351276 590730 351876 6 vssa1
port 535 nsew ground input
rlabel metal5 s -6806 387276 590730 387876 6 vssa1
port 535 nsew ground input
rlabel metal5 s -6806 423276 590730 423876 6 vssa1
port 535 nsew ground input
rlabel metal5 s -6806 459276 590730 459876 6 vssa1
port 535 nsew ground input
rlabel metal5 s -6806 495276 590730 495876 6 vssa1
port 535 nsew ground input
rlabel metal5 s -6806 531276 590730 531876 6 vssa1
port 535 nsew ground input
rlabel metal5 s -6806 567276 590730 567876 6 vssa1
port 535 nsew ground input
rlabel metal5 s -6806 603276 590730 603876 6 vssa1
port 535 nsew ground input
rlabel metal5 s -6806 639276 590730 639876 6 vssa1
port 535 nsew ground input
rlabel metal5 s -6806 675276 590730 675876 6 vssa1
port 535 nsew ground input
rlabel metal5 s -6806 709050 590730 709670 6 vssa1
port 535 nsew ground input
rlabel metal4 s 62204 -5734 62804 38000 6 vssa1
port 535 nsew ground input
rlabel metal4 s 98204 -5734 98804 38000 6 vssa1
port 535 nsew ground input
rlabel metal4 s 134204 -5734 134804 38000 6 vssa1
port 535 nsew ground input
rlabel metal4 s 170204 -5734 170804 38000 6 vssa1
port 535 nsew ground input
rlabel metal4 s 206204 -5734 206804 38000 6 vssa1
port 535 nsew ground input
rlabel metal4 s 62204 242304 62804 338000 6 vssa1
port 535 nsew ground input
rlabel metal4 s 98204 242304 98804 338000 6 vssa1
port 535 nsew ground input
rlabel metal4 s 134204 242304 134804 338000 6 vssa1
port 535 nsew ground input
rlabel metal4 s 170204 242304 170804 338000 6 vssa1
port 535 nsew ground input
rlabel metal4 s 350204 -5734 350804 338000 6 vssa1
port 535 nsew ground input
rlabel metal4 s 386204 -5734 386804 338000 6 vssa1
port 535 nsew ground input
rlabel metal4 s 422204 -5734 422804 338000 6 vssa1
port 535 nsew ground input
rlabel metal4 s 458204 -5734 458804 338000 6 vssa1
port 535 nsew ground input
rlabel metal4 s -6806 -5734 -6186 709670 4 vssa1
port 535 nsew ground input
rlabel metal4 s 26204 -5734 26804 709670 6 vssa1
port 535 nsew ground input
rlabel metal4 s 62204 425308 62804 709670 6 vssa1
port 535 nsew ground input
rlabel metal4 s 98204 425308 98804 709670 6 vssa1
port 535 nsew ground input
rlabel metal4 s 134204 425308 134804 709670 6 vssa1
port 535 nsew ground input
rlabel metal4 s 170204 425308 170804 709670 6 vssa1
port 535 nsew ground input
rlabel metal4 s 206204 242304 206804 709670 6 vssa1
port 535 nsew ground input
rlabel metal4 s 242204 -5734 242804 709670 6 vssa1
port 535 nsew ground input
rlabel metal4 s 278204 -5734 278804 709670 6 vssa1
port 535 nsew ground input
rlabel metal4 s 314204 -5734 314804 709670 6 vssa1
port 535 nsew ground input
rlabel metal4 s 350204 425308 350804 709670 6 vssa1
port 535 nsew ground input
rlabel metal4 s 386204 425308 386804 709670 6 vssa1
port 535 nsew ground input
rlabel metal4 s 422204 425308 422804 709670 6 vssa1
port 535 nsew ground input
rlabel metal4 s 458204 425308 458804 709670 6 vssa1
port 535 nsew ground input
rlabel metal4 s 494204 -5734 494804 709670 6 vssa1
port 535 nsew ground input
rlabel metal4 s 530204 -5734 530804 709670 6 vssa1
port 535 nsew ground input
rlabel metal4 s 566204 -5734 566804 709670 6 vssa1
port 535 nsew ground input
rlabel metal4 s 590110 -5734 590730 709670 6 vssa1
port 535 nsew ground input
rlabel metal5 s -8726 -7654 592650 -7034 8 vssa2
port 536 nsew ground input
rlabel metal5 s -8726 30976 592650 31576 6 vssa2
port 536 nsew ground input
rlabel metal5 s -8726 66976 592650 67576 6 vssa2
port 536 nsew ground input
rlabel metal5 s -8726 102976 592650 103576 6 vssa2
port 536 nsew ground input
rlabel metal5 s -8726 138976 592650 139576 6 vssa2
port 536 nsew ground input
rlabel metal5 s -8726 174976 592650 175576 6 vssa2
port 536 nsew ground input
rlabel metal5 s -8726 210976 592650 211576 6 vssa2
port 536 nsew ground input
rlabel metal5 s -8726 246976 592650 247576 6 vssa2
port 536 nsew ground input
rlabel metal5 s -8726 282976 592650 283576 6 vssa2
port 536 nsew ground input
rlabel metal5 s -8726 318976 592650 319576 6 vssa2
port 536 nsew ground input
rlabel metal5 s -8726 354976 592650 355576 6 vssa2
port 536 nsew ground input
rlabel metal5 s -8726 390976 592650 391576 6 vssa2
port 536 nsew ground input
rlabel metal5 s -8726 426976 592650 427576 6 vssa2
port 536 nsew ground input
rlabel metal5 s -8726 462976 592650 463576 6 vssa2
port 536 nsew ground input
rlabel metal5 s -8726 498976 592650 499576 6 vssa2
port 536 nsew ground input
rlabel metal5 s -8726 534976 592650 535576 6 vssa2
port 536 nsew ground input
rlabel metal5 s -8726 570976 592650 571576 6 vssa2
port 536 nsew ground input
rlabel metal5 s -8726 606976 592650 607576 6 vssa2
port 536 nsew ground input
rlabel metal5 s -8726 642976 592650 643576 6 vssa2
port 536 nsew ground input
rlabel metal5 s -8726 678976 592650 679576 6 vssa2
port 536 nsew ground input
rlabel metal5 s -8726 710970 592650 711590 6 vssa2
port 536 nsew ground input
rlabel metal4 s 65904 -7654 66504 38000 6 vssa2
port 536 nsew ground input
rlabel metal4 s 101904 -7654 102504 38000 6 vssa2
port 536 nsew ground input
rlabel metal4 s 137904 -7654 138504 38000 6 vssa2
port 536 nsew ground input
rlabel metal4 s 173904 -7654 174504 38000 6 vssa2
port 536 nsew ground input
rlabel metal4 s 209904 -7654 210504 38000 6 vssa2
port 536 nsew ground input
rlabel metal4 s 65904 242304 66504 338000 6 vssa2
port 536 nsew ground input
rlabel metal4 s 101904 242304 102504 338000 6 vssa2
port 536 nsew ground input
rlabel metal4 s 137904 242304 138504 338000 6 vssa2
port 536 nsew ground input
rlabel metal4 s 173904 242304 174504 338000 6 vssa2
port 536 nsew ground input
rlabel metal4 s 353904 -7654 354504 338000 6 vssa2
port 536 nsew ground input
rlabel metal4 s 389904 -7654 390504 338000 6 vssa2
port 536 nsew ground input
rlabel metal4 s 425904 -7654 426504 338000 6 vssa2
port 536 nsew ground input
rlabel metal4 s 461904 -7654 462504 338000 6 vssa2
port 536 nsew ground input
rlabel metal4 s -8726 -7654 -8106 711590 4 vssa2
port 536 nsew ground input
rlabel metal4 s 29904 -7654 30504 711590 6 vssa2
port 536 nsew ground input
rlabel metal4 s 65904 425308 66504 711590 6 vssa2
port 536 nsew ground input
rlabel metal4 s 101904 425308 102504 711590 6 vssa2
port 536 nsew ground input
rlabel metal4 s 137904 425308 138504 711590 6 vssa2
port 536 nsew ground input
rlabel metal4 s 173904 425308 174504 711590 6 vssa2
port 536 nsew ground input
rlabel metal4 s 209904 242304 210504 711590 6 vssa2
port 536 nsew ground input
rlabel metal4 s 245904 -7654 246504 711590 6 vssa2
port 536 nsew ground input
rlabel metal4 s 281904 -7654 282504 711590 6 vssa2
port 536 nsew ground input
rlabel metal4 s 317904 -7654 318504 711590 6 vssa2
port 536 nsew ground input
rlabel metal4 s 353904 425308 354504 711590 6 vssa2
port 536 nsew ground input
rlabel metal4 s 389904 425308 390504 711590 6 vssa2
port 536 nsew ground input
rlabel metal4 s 425904 425308 426504 711590 6 vssa2
port 536 nsew ground input
rlabel metal4 s 461904 425308 462504 711590 6 vssa2
port 536 nsew ground input
rlabel metal4 s 497904 -7654 498504 711590 6 vssa2
port 536 nsew ground input
rlabel metal4 s 533904 -7654 534504 711590 6 vssa2
port 536 nsew ground input
rlabel metal4 s 569904 -7654 570504 711590 6 vssa2
port 536 nsew ground input
rlabel metal4 s 592030 -7654 592650 711590 6 vssa2
port 536 nsew ground input
rlabel metal5 s -2966 -1894 586890 -1274 8 vssd1
port 537 nsew ground input
rlabel metal5 s -2966 19876 586890 20476 6 vssd1
port 537 nsew ground input
rlabel metal5 s -2966 55876 586890 56476 6 vssd1
port 537 nsew ground input
rlabel metal5 s -2966 91876 586890 92476 6 vssd1
port 537 nsew ground input
rlabel metal5 s -2966 127876 586890 128476 6 vssd1
port 537 nsew ground input
rlabel metal5 s -2966 163876 586890 164476 6 vssd1
port 537 nsew ground input
rlabel metal5 s -2966 199876 586890 200476 6 vssd1
port 537 nsew ground input
rlabel metal5 s -2966 235876 586890 236476 6 vssd1
port 537 nsew ground input
rlabel metal5 s -2966 271876 586890 272476 6 vssd1
port 537 nsew ground input
rlabel metal5 s -2966 307876 586890 308476 6 vssd1
port 537 nsew ground input
rlabel metal5 s -2966 343876 586890 344476 6 vssd1
port 537 nsew ground input
rlabel metal5 s -2966 379876 586890 380476 6 vssd1
port 537 nsew ground input
rlabel metal5 s -2966 415876 586890 416476 6 vssd1
port 537 nsew ground input
rlabel metal5 s -2966 451876 586890 452476 6 vssd1
port 537 nsew ground input
rlabel metal5 s -2966 487876 586890 488476 6 vssd1
port 537 nsew ground input
rlabel metal5 s -2966 523876 586890 524476 6 vssd1
port 537 nsew ground input
rlabel metal5 s -2966 559876 586890 560476 6 vssd1
port 537 nsew ground input
rlabel metal5 s -2966 595876 586890 596476 6 vssd1
port 537 nsew ground input
rlabel metal5 s -2966 631876 586890 632476 6 vssd1
port 537 nsew ground input
rlabel metal5 s -2966 667876 586890 668476 6 vssd1
port 537 nsew ground input
rlabel metal5 s -2966 705210 586890 705830 6 vssd1
port 537 nsew ground input
rlabel metal4 s 54804 -1894 55404 38000 6 vssd1
port 537 nsew ground input
rlabel metal4 s 90804 -1894 91404 38000 6 vssd1
port 537 nsew ground input
rlabel metal4 s 126804 -1894 127404 38000 6 vssd1
port 537 nsew ground input
rlabel metal4 s 162804 -1894 163404 38000 6 vssd1
port 537 nsew ground input
rlabel metal4 s 198804 -1894 199404 38000 6 vssd1
port 537 nsew ground input
rlabel metal4 s 234804 -1894 235404 38000 6 vssd1
port 537 nsew ground input
rlabel metal4 s 54804 242304 55404 338000 6 vssd1
port 537 nsew ground input
rlabel metal4 s 90804 242304 91404 338000 6 vssd1
port 537 nsew ground input
rlabel metal4 s 126804 242304 127404 338000 6 vssd1
port 537 nsew ground input
rlabel metal4 s 162804 242304 163404 338000 6 vssd1
port 537 nsew ground input
rlabel metal4 s 342804 -1894 343404 338000 6 vssd1
port 537 nsew ground input
rlabel metal4 s 378804 -1894 379404 338000 6 vssd1
port 537 nsew ground input
rlabel metal4 s 414804 -1894 415404 338000 6 vssd1
port 537 nsew ground input
rlabel metal4 s 450804 -1894 451404 338000 6 vssd1
port 537 nsew ground input
rlabel metal4 s -2966 -1894 -2346 705830 4 vssd1
port 537 nsew ground input
rlabel metal4 s 18804 -1894 19404 705830 6 vssd1
port 537 nsew ground input
rlabel metal4 s 54804 425308 55404 705830 6 vssd1
port 537 nsew ground input
rlabel metal4 s 90804 425308 91404 705830 6 vssd1
port 537 nsew ground input
rlabel metal4 s 126804 425308 127404 705830 6 vssd1
port 537 nsew ground input
rlabel metal4 s 162804 425308 163404 705830 6 vssd1
port 537 nsew ground input
rlabel metal4 s 198804 242304 199404 705830 6 vssd1
port 537 nsew ground input
rlabel metal4 s 234804 242304 235404 705830 6 vssd1
port 537 nsew ground input
rlabel metal4 s 270804 -1894 271404 705830 6 vssd1
port 537 nsew ground input
rlabel metal4 s 306804 -1894 307404 705830 6 vssd1
port 537 nsew ground input
rlabel metal4 s 342804 425308 343404 705830 6 vssd1
port 537 nsew ground input
rlabel metal4 s 378804 425308 379404 705830 6 vssd1
port 537 nsew ground input
rlabel metal4 s 414804 425308 415404 705830 6 vssd1
port 537 nsew ground input
rlabel metal4 s 450804 425308 451404 705830 6 vssd1
port 537 nsew ground input
rlabel metal4 s 486804 -1894 487404 705830 6 vssd1
port 537 nsew ground input
rlabel metal4 s 522804 -1894 523404 705830 6 vssd1
port 537 nsew ground input
rlabel metal4 s 558804 -1894 559404 705830 6 vssd1
port 537 nsew ground input
rlabel metal4 s 586270 -1894 586890 705830 6 vssd1
port 537 nsew ground input
rlabel metal5 s -4886 -3814 588810 -3194 8 vssd2
port 538 nsew ground input
rlabel metal5 s -4886 23576 588810 24176 6 vssd2
port 538 nsew ground input
rlabel metal5 s -4886 59576 588810 60176 6 vssd2
port 538 nsew ground input
rlabel metal5 s -4886 95576 588810 96176 6 vssd2
port 538 nsew ground input
rlabel metal5 s -4886 131576 588810 132176 6 vssd2
port 538 nsew ground input
rlabel metal5 s -4886 167576 588810 168176 6 vssd2
port 538 nsew ground input
rlabel metal5 s -4886 203576 588810 204176 6 vssd2
port 538 nsew ground input
rlabel metal5 s -4886 239576 588810 240176 6 vssd2
port 538 nsew ground input
rlabel metal5 s -4886 275576 588810 276176 6 vssd2
port 538 nsew ground input
rlabel metal5 s -4886 311576 588810 312176 6 vssd2
port 538 nsew ground input
rlabel metal5 s -4886 347576 588810 348176 6 vssd2
port 538 nsew ground input
rlabel metal5 s -4886 383576 588810 384176 6 vssd2
port 538 nsew ground input
rlabel metal5 s -4886 419576 588810 420176 6 vssd2
port 538 nsew ground input
rlabel metal5 s -4886 455576 588810 456176 6 vssd2
port 538 nsew ground input
rlabel metal5 s -4886 491576 588810 492176 6 vssd2
port 538 nsew ground input
rlabel metal5 s -4886 527576 588810 528176 6 vssd2
port 538 nsew ground input
rlabel metal5 s -4886 563576 588810 564176 6 vssd2
port 538 nsew ground input
rlabel metal5 s -4886 599576 588810 600176 6 vssd2
port 538 nsew ground input
rlabel metal5 s -4886 635576 588810 636176 6 vssd2
port 538 nsew ground input
rlabel metal5 s -4886 671576 588810 672176 6 vssd2
port 538 nsew ground input
rlabel metal5 s -4886 707130 588810 707750 6 vssd2
port 538 nsew ground input
rlabel metal4 s 58504 -3814 59104 38000 6 vssd2
port 538 nsew ground input
rlabel metal4 s 94504 -3814 95104 38000 6 vssd2
port 538 nsew ground input
rlabel metal4 s 130504 -3814 131104 38000 6 vssd2
port 538 nsew ground input
rlabel metal4 s 166504 -3814 167104 38000 6 vssd2
port 538 nsew ground input
rlabel metal4 s 202504 -3814 203104 38000 6 vssd2
port 538 nsew ground input
rlabel metal4 s 238504 -3814 239104 38000 6 vssd2
port 538 nsew ground input
rlabel metal4 s 58504 242304 59104 338000 6 vssd2
port 538 nsew ground input
rlabel metal4 s 94504 242304 95104 338000 6 vssd2
port 538 nsew ground input
rlabel metal4 s 130504 242304 131104 338000 6 vssd2
port 538 nsew ground input
rlabel metal4 s 166504 242304 167104 338000 6 vssd2
port 538 nsew ground input
rlabel metal4 s 346504 -3814 347104 338000 6 vssd2
port 538 nsew ground input
rlabel metal4 s 382504 -3814 383104 338000 6 vssd2
port 538 nsew ground input
rlabel metal4 s 418504 -3814 419104 338000 6 vssd2
port 538 nsew ground input
rlabel metal4 s 454504 -3814 455104 338000 6 vssd2
port 538 nsew ground input
rlabel metal4 s -4886 -3814 -4266 707750 4 vssd2
port 538 nsew ground input
rlabel metal4 s 22504 -3814 23104 707750 6 vssd2
port 538 nsew ground input
rlabel metal4 s 58504 425308 59104 707750 6 vssd2
port 538 nsew ground input
rlabel metal4 s 94504 425308 95104 707750 6 vssd2
port 538 nsew ground input
rlabel metal4 s 130504 425308 131104 707750 6 vssd2
port 538 nsew ground input
rlabel metal4 s 166504 425308 167104 707750 6 vssd2
port 538 nsew ground input
rlabel metal4 s 202504 242304 203104 707750 6 vssd2
port 538 nsew ground input
rlabel metal4 s 238504 242304 239104 707750 6 vssd2
port 538 nsew ground input
rlabel metal4 s 274504 -3814 275104 707750 6 vssd2
port 538 nsew ground input
rlabel metal4 s 310504 -3814 311104 707750 6 vssd2
port 538 nsew ground input
rlabel metal4 s 346504 425308 347104 707750 6 vssd2
port 538 nsew ground input
rlabel metal4 s 382504 425308 383104 707750 6 vssd2
port 538 nsew ground input
rlabel metal4 s 418504 425308 419104 707750 6 vssd2
port 538 nsew ground input
rlabel metal4 s 454504 425308 455104 707750 6 vssd2
port 538 nsew ground input
rlabel metal4 s 490504 -3814 491104 707750 6 vssd2
port 538 nsew ground input
rlabel metal4 s 526504 -3814 527104 707750 6 vssd2
port 538 nsew ground input
rlabel metal4 s 562504 -3814 563104 707750 6 vssd2
port 538 nsew ground input
rlabel metal4 s 588190 -3814 588810 707750 6 vssd2
port 538 nsew ground input
rlabel metal2 s 542 -960 654 480 8 wb_clk_i
port 539 nsew signal input
rlabel metal2 s 1646 -960 1758 480 8 wb_rst_i
port 540 nsew signal input
rlabel metal2 s 2842 -960 2954 480 8 wbs_ack_o
port 541 nsew signal tristate
rlabel metal2 s 7626 -960 7738 480 8 wbs_adr_i[0]
port 542 nsew signal input
rlabel metal2 s 47830 -960 47942 480 8 wbs_adr_i[10]
port 543 nsew signal input
rlabel metal2 s 51326 -960 51438 480 8 wbs_adr_i[11]
port 544 nsew signal input
rlabel metal2 s 54914 -960 55026 480 8 wbs_adr_i[12]
port 545 nsew signal input
rlabel metal2 s 58410 -960 58522 480 8 wbs_adr_i[13]
port 546 nsew signal input
rlabel metal2 s 61998 -960 62110 480 8 wbs_adr_i[14]
port 547 nsew signal input
rlabel metal2 s 65494 -960 65606 480 8 wbs_adr_i[15]
port 548 nsew signal input
rlabel metal2 s 69082 -960 69194 480 8 wbs_adr_i[16]
port 549 nsew signal input
rlabel metal2 s 72578 -960 72690 480 8 wbs_adr_i[17]
port 550 nsew signal input
rlabel metal2 s 76166 -960 76278 480 8 wbs_adr_i[18]
port 551 nsew signal input
rlabel metal2 s 79662 -960 79774 480 8 wbs_adr_i[19]
port 552 nsew signal input
rlabel metal2 s 12318 -960 12430 480 8 wbs_adr_i[1]
port 553 nsew signal input
rlabel metal2 s 83250 -960 83362 480 8 wbs_adr_i[20]
port 554 nsew signal input
rlabel metal2 s 86838 -960 86950 480 8 wbs_adr_i[21]
port 555 nsew signal input
rlabel metal2 s 90334 -960 90446 480 8 wbs_adr_i[22]
port 556 nsew signal input
rlabel metal2 s 93922 -960 94034 480 8 wbs_adr_i[23]
port 557 nsew signal input
rlabel metal2 s 97418 -960 97530 480 8 wbs_adr_i[24]
port 558 nsew signal input
rlabel metal2 s 101006 -960 101118 480 8 wbs_adr_i[25]
port 559 nsew signal input
rlabel metal2 s 104502 -960 104614 480 8 wbs_adr_i[26]
port 560 nsew signal input
rlabel metal2 s 108090 -960 108202 480 8 wbs_adr_i[27]
port 561 nsew signal input
rlabel metal2 s 111586 -960 111698 480 8 wbs_adr_i[28]
port 562 nsew signal input
rlabel metal2 s 115174 -960 115286 480 8 wbs_adr_i[29]
port 563 nsew signal input
rlabel metal2 s 17010 -960 17122 480 8 wbs_adr_i[2]
port 564 nsew signal input
rlabel metal2 s 118762 -960 118874 480 8 wbs_adr_i[30]
port 565 nsew signal input
rlabel metal2 s 122258 -960 122370 480 8 wbs_adr_i[31]
port 566 nsew signal input
rlabel metal2 s 21794 -960 21906 480 8 wbs_adr_i[3]
port 567 nsew signal input
rlabel metal2 s 26486 -960 26598 480 8 wbs_adr_i[4]
port 568 nsew signal input
rlabel metal2 s 30074 -960 30186 480 8 wbs_adr_i[5]
port 569 nsew signal input
rlabel metal2 s 33570 -960 33682 480 8 wbs_adr_i[6]
port 570 nsew signal input
rlabel metal2 s 37158 -960 37270 480 8 wbs_adr_i[7]
port 571 nsew signal input
rlabel metal2 s 40654 -960 40766 480 8 wbs_adr_i[8]
port 572 nsew signal input
rlabel metal2 s 44242 -960 44354 480 8 wbs_adr_i[9]
port 573 nsew signal input
rlabel metal2 s 4038 -960 4150 480 8 wbs_cyc_i
port 574 nsew signal input
rlabel metal2 s 8730 -960 8842 480 8 wbs_dat_i[0]
port 575 nsew signal input
rlabel metal2 s 48934 -960 49046 480 8 wbs_dat_i[10]
port 576 nsew signal input
rlabel metal2 s 52522 -960 52634 480 8 wbs_dat_i[11]
port 577 nsew signal input
rlabel metal2 s 56018 -960 56130 480 8 wbs_dat_i[12]
port 578 nsew signal input
rlabel metal2 s 59606 -960 59718 480 8 wbs_dat_i[13]
port 579 nsew signal input
rlabel metal2 s 63194 -960 63306 480 8 wbs_dat_i[14]
port 580 nsew signal input
rlabel metal2 s 66690 -960 66802 480 8 wbs_dat_i[15]
port 581 nsew signal input
rlabel metal2 s 70278 -960 70390 480 8 wbs_dat_i[16]
port 582 nsew signal input
rlabel metal2 s 73774 -960 73886 480 8 wbs_dat_i[17]
port 583 nsew signal input
rlabel metal2 s 77362 -960 77474 480 8 wbs_dat_i[18]
port 584 nsew signal input
rlabel metal2 s 80858 -960 80970 480 8 wbs_dat_i[19]
port 585 nsew signal input
rlabel metal2 s 13514 -960 13626 480 8 wbs_dat_i[1]
port 586 nsew signal input
rlabel metal2 s 84446 -960 84558 480 8 wbs_dat_i[20]
port 587 nsew signal input
rlabel metal2 s 87942 -960 88054 480 8 wbs_dat_i[21]
port 588 nsew signal input
rlabel metal2 s 91530 -960 91642 480 8 wbs_dat_i[22]
port 589 nsew signal input
rlabel metal2 s 95118 -960 95230 480 8 wbs_dat_i[23]
port 590 nsew signal input
rlabel metal2 s 98614 -960 98726 480 8 wbs_dat_i[24]
port 591 nsew signal input
rlabel metal2 s 102202 -960 102314 480 8 wbs_dat_i[25]
port 592 nsew signal input
rlabel metal2 s 105698 -960 105810 480 8 wbs_dat_i[26]
port 593 nsew signal input
rlabel metal2 s 109286 -960 109398 480 8 wbs_dat_i[27]
port 594 nsew signal input
rlabel metal2 s 112782 -960 112894 480 8 wbs_dat_i[28]
port 595 nsew signal input
rlabel metal2 s 116370 -960 116482 480 8 wbs_dat_i[29]
port 596 nsew signal input
rlabel metal2 s 18206 -960 18318 480 8 wbs_dat_i[2]
port 597 nsew signal input
rlabel metal2 s 119866 -960 119978 480 8 wbs_dat_i[30]
port 598 nsew signal input
rlabel metal2 s 123454 -960 123566 480 8 wbs_dat_i[31]
port 599 nsew signal input
rlabel metal2 s 22990 -960 23102 480 8 wbs_dat_i[3]
port 600 nsew signal input
rlabel metal2 s 27682 -960 27794 480 8 wbs_dat_i[4]
port 601 nsew signal input
rlabel metal2 s 31270 -960 31382 480 8 wbs_dat_i[5]
port 602 nsew signal input
rlabel metal2 s 34766 -960 34878 480 8 wbs_dat_i[6]
port 603 nsew signal input
rlabel metal2 s 38354 -960 38466 480 8 wbs_dat_i[7]
port 604 nsew signal input
rlabel metal2 s 41850 -960 41962 480 8 wbs_dat_i[8]
port 605 nsew signal input
rlabel metal2 s 45438 -960 45550 480 8 wbs_dat_i[9]
port 606 nsew signal input
rlabel metal2 s 9926 -960 10038 480 8 wbs_dat_o[0]
port 607 nsew signal tristate
rlabel metal2 s 50130 -960 50242 480 8 wbs_dat_o[10]
port 608 nsew signal tristate
rlabel metal2 s 53718 -960 53830 480 8 wbs_dat_o[11]
port 609 nsew signal tristate
rlabel metal2 s 57214 -960 57326 480 8 wbs_dat_o[12]
port 610 nsew signal tristate
rlabel metal2 s 60802 -960 60914 480 8 wbs_dat_o[13]
port 611 nsew signal tristate
rlabel metal2 s 64298 -960 64410 480 8 wbs_dat_o[14]
port 612 nsew signal tristate
rlabel metal2 s 67886 -960 67998 480 8 wbs_dat_o[15]
port 613 nsew signal tristate
rlabel metal2 s 71474 -960 71586 480 8 wbs_dat_o[16]
port 614 nsew signal tristate
rlabel metal2 s 74970 -960 75082 480 8 wbs_dat_o[17]
port 615 nsew signal tristate
rlabel metal2 s 78558 -960 78670 480 8 wbs_dat_o[18]
port 616 nsew signal tristate
rlabel metal2 s 82054 -960 82166 480 8 wbs_dat_o[19]
port 617 nsew signal tristate
rlabel metal2 s 14710 -960 14822 480 8 wbs_dat_o[1]
port 618 nsew signal tristate
rlabel metal2 s 85642 -960 85754 480 8 wbs_dat_o[20]
port 619 nsew signal tristate
rlabel metal2 s 89138 -960 89250 480 8 wbs_dat_o[21]
port 620 nsew signal tristate
rlabel metal2 s 92726 -960 92838 480 8 wbs_dat_o[22]
port 621 nsew signal tristate
rlabel metal2 s 96222 -960 96334 480 8 wbs_dat_o[23]
port 622 nsew signal tristate
rlabel metal2 s 99810 -960 99922 480 8 wbs_dat_o[24]
port 623 nsew signal tristate
rlabel metal2 s 103306 -960 103418 480 8 wbs_dat_o[25]
port 624 nsew signal tristate
rlabel metal2 s 106894 -960 107006 480 8 wbs_dat_o[26]
port 625 nsew signal tristate
rlabel metal2 s 110482 -960 110594 480 8 wbs_dat_o[27]
port 626 nsew signal tristate
rlabel metal2 s 113978 -960 114090 480 8 wbs_dat_o[28]
port 627 nsew signal tristate
rlabel metal2 s 117566 -960 117678 480 8 wbs_dat_o[29]
port 628 nsew signal tristate
rlabel metal2 s 19402 -960 19514 480 8 wbs_dat_o[2]
port 629 nsew signal tristate
rlabel metal2 s 121062 -960 121174 480 8 wbs_dat_o[30]
port 630 nsew signal tristate
rlabel metal2 s 124650 -960 124762 480 8 wbs_dat_o[31]
port 631 nsew signal tristate
rlabel metal2 s 24186 -960 24298 480 8 wbs_dat_o[3]
port 632 nsew signal tristate
rlabel metal2 s 28878 -960 28990 480 8 wbs_dat_o[4]
port 633 nsew signal tristate
rlabel metal2 s 32374 -960 32486 480 8 wbs_dat_o[5]
port 634 nsew signal tristate
rlabel metal2 s 35962 -960 36074 480 8 wbs_dat_o[6]
port 635 nsew signal tristate
rlabel metal2 s 39550 -960 39662 480 8 wbs_dat_o[7]
port 636 nsew signal tristate
rlabel metal2 s 43046 -960 43158 480 8 wbs_dat_o[8]
port 637 nsew signal tristate
rlabel metal2 s 46634 -960 46746 480 8 wbs_dat_o[9]
port 638 nsew signal tristate
rlabel metal2 s 11122 -960 11234 480 8 wbs_sel_i[0]
port 639 nsew signal input
rlabel metal2 s 15906 -960 16018 480 8 wbs_sel_i[1]
port 640 nsew signal input
rlabel metal2 s 20598 -960 20710 480 8 wbs_sel_i[2]
port 641 nsew signal input
rlabel metal2 s 25290 -960 25402 480 8 wbs_sel_i[3]
port 642 nsew signal input
rlabel metal2 s 5234 -960 5346 480 8 wbs_stb_i
port 643 nsew signal input
rlabel metal2 s 6430 -960 6542 480 8 wbs_we_i
port 644 nsew signal input
<< properties >>
string FIXED_BBOX 0 0 584000 704000
<< end >>
