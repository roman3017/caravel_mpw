magic
tech sky130A
magscale 1 2
timestamp 1645327450
<< obsli1 >>
rect 1104 2159 197955 198033
<< obsm1 >>
rect 1026 348 197967 198064
<< metal2 >>
rect 570 199504 626 200304
rect 1766 199504 1822 200304
rect 3054 199504 3110 200304
rect 4342 199504 4398 200304
rect 5630 199504 5686 200304
rect 6918 199504 6974 200304
rect 8206 199504 8262 200304
rect 9494 199504 9550 200304
rect 10782 199504 10838 200304
rect 12070 199504 12126 200304
rect 13266 199504 13322 200304
rect 14554 199504 14610 200304
rect 15842 199504 15898 200304
rect 17130 199504 17186 200304
rect 18418 199504 18474 200304
rect 19706 199504 19762 200304
rect 20994 199504 21050 200304
rect 22282 199504 22338 200304
rect 23570 199504 23626 200304
rect 24858 199504 24914 200304
rect 26054 199504 26110 200304
rect 27342 199504 27398 200304
rect 28630 199504 28686 200304
rect 29918 199504 29974 200304
rect 31206 199504 31262 200304
rect 32494 199504 32550 200304
rect 33782 199504 33838 200304
rect 35070 199504 35126 200304
rect 36358 199504 36414 200304
rect 37646 199504 37702 200304
rect 38842 199504 38898 200304
rect 40130 199504 40186 200304
rect 41418 199504 41474 200304
rect 42706 199504 42762 200304
rect 43994 199504 44050 200304
rect 45282 199504 45338 200304
rect 46570 199504 46626 200304
rect 47858 199504 47914 200304
rect 49146 199504 49202 200304
rect 50342 199504 50398 200304
rect 51630 199504 51686 200304
rect 52918 199504 52974 200304
rect 54206 199504 54262 200304
rect 55494 199504 55550 200304
rect 56782 199504 56838 200304
rect 58070 199504 58126 200304
rect 59358 199504 59414 200304
rect 60646 199504 60702 200304
rect 61934 199504 61990 200304
rect 63130 199504 63186 200304
rect 64418 199504 64474 200304
rect 65706 199504 65762 200304
rect 66994 199504 67050 200304
rect 68282 199504 68338 200304
rect 69570 199504 69626 200304
rect 70858 199504 70914 200304
rect 72146 199504 72202 200304
rect 73434 199504 73490 200304
rect 74722 199504 74778 200304
rect 75918 199504 75974 200304
rect 77206 199504 77262 200304
rect 78494 199504 78550 200304
rect 79782 199504 79838 200304
rect 81070 199504 81126 200304
rect 82358 199504 82414 200304
rect 83646 199504 83702 200304
rect 84934 199504 84990 200304
rect 86222 199504 86278 200304
rect 87418 199504 87474 200304
rect 88706 199504 88762 200304
rect 89994 199504 90050 200304
rect 91282 199504 91338 200304
rect 92570 199504 92626 200304
rect 93858 199504 93914 200304
rect 95146 199504 95202 200304
rect 96434 199504 96490 200304
rect 97722 199504 97778 200304
rect 99010 199504 99066 200304
rect 100206 199504 100262 200304
rect 101494 199504 101550 200304
rect 102782 199504 102838 200304
rect 104070 199504 104126 200304
rect 105358 199504 105414 200304
rect 106646 199504 106702 200304
rect 107934 199504 107990 200304
rect 109222 199504 109278 200304
rect 110510 199504 110566 200304
rect 111798 199504 111854 200304
rect 112994 199504 113050 200304
rect 114282 199504 114338 200304
rect 115570 199504 115626 200304
rect 116858 199504 116914 200304
rect 118146 199504 118202 200304
rect 119434 199504 119490 200304
rect 120722 199504 120778 200304
rect 122010 199504 122066 200304
rect 123298 199504 123354 200304
rect 124494 199504 124550 200304
rect 125782 199504 125838 200304
rect 127070 199504 127126 200304
rect 128358 199504 128414 200304
rect 129646 199504 129702 200304
rect 130934 199504 130990 200304
rect 132222 199504 132278 200304
rect 133510 199504 133566 200304
rect 134798 199504 134854 200304
rect 136086 199504 136142 200304
rect 137282 199504 137338 200304
rect 138570 199504 138626 200304
rect 139858 199504 139914 200304
rect 141146 199504 141202 200304
rect 142434 199504 142490 200304
rect 143722 199504 143778 200304
rect 145010 199504 145066 200304
rect 146298 199504 146354 200304
rect 147586 199504 147642 200304
rect 148874 199504 148930 200304
rect 150070 199504 150126 200304
rect 151358 199504 151414 200304
rect 152646 199504 152702 200304
rect 153934 199504 153990 200304
rect 155222 199504 155278 200304
rect 156510 199504 156566 200304
rect 157798 199504 157854 200304
rect 159086 199504 159142 200304
rect 160374 199504 160430 200304
rect 161570 199504 161626 200304
rect 162858 199504 162914 200304
rect 164146 199504 164202 200304
rect 165434 199504 165490 200304
rect 166722 199504 166778 200304
rect 168010 199504 168066 200304
rect 169298 199504 169354 200304
rect 170586 199504 170642 200304
rect 171874 199504 171930 200304
rect 173162 199504 173218 200304
rect 174358 199504 174414 200304
rect 175646 199504 175702 200304
rect 176934 199504 176990 200304
rect 178222 199504 178278 200304
rect 179510 199504 179566 200304
rect 180798 199504 180854 200304
rect 182086 199504 182142 200304
rect 183374 199504 183430 200304
rect 184662 199504 184718 200304
rect 185950 199504 186006 200304
rect 187146 199504 187202 200304
rect 188434 199504 188490 200304
rect 189722 199504 189778 200304
rect 191010 199504 191066 200304
rect 192298 199504 192354 200304
rect 193586 199504 193642 200304
rect 194874 199504 194930 200304
rect 196162 199504 196218 200304
rect 197450 199504 197506 200304
rect 662 0 718 800
rect 1950 0 2006 800
rect 3238 0 3294 800
rect 4526 0 4582 800
rect 5906 0 5962 800
rect 7194 0 7250 800
rect 8482 0 8538 800
rect 9770 0 9826 800
rect 11150 0 11206 800
rect 12438 0 12494 800
rect 13726 0 13782 800
rect 15014 0 15070 800
rect 16394 0 16450 800
rect 17682 0 17738 800
rect 18970 0 19026 800
rect 20258 0 20314 800
rect 21638 0 21694 800
rect 22926 0 22982 800
rect 24214 0 24270 800
rect 25594 0 25650 800
rect 26882 0 26938 800
rect 28170 0 28226 800
rect 29458 0 29514 800
rect 30838 0 30894 800
rect 32126 0 32182 800
rect 33414 0 33470 800
rect 34702 0 34758 800
rect 36082 0 36138 800
rect 37370 0 37426 800
rect 38658 0 38714 800
rect 39946 0 40002 800
rect 41326 0 41382 800
rect 42614 0 42670 800
rect 43902 0 43958 800
rect 45282 0 45338 800
rect 46570 0 46626 800
rect 47858 0 47914 800
rect 49146 0 49202 800
rect 50526 0 50582 800
rect 51814 0 51870 800
rect 53102 0 53158 800
rect 54390 0 54446 800
rect 55770 0 55826 800
rect 57058 0 57114 800
rect 58346 0 58402 800
rect 59634 0 59690 800
rect 61014 0 61070 800
rect 62302 0 62358 800
rect 63590 0 63646 800
rect 64878 0 64934 800
rect 66258 0 66314 800
rect 67546 0 67602 800
rect 68834 0 68890 800
rect 70214 0 70270 800
rect 71502 0 71558 800
rect 72790 0 72846 800
rect 74078 0 74134 800
rect 75458 0 75514 800
rect 76746 0 76802 800
rect 78034 0 78090 800
rect 79322 0 79378 800
rect 80702 0 80758 800
rect 81990 0 82046 800
rect 83278 0 83334 800
rect 84566 0 84622 800
rect 85946 0 86002 800
rect 87234 0 87290 800
rect 88522 0 88578 800
rect 89902 0 89958 800
rect 91190 0 91246 800
rect 92478 0 92534 800
rect 93766 0 93822 800
rect 95146 0 95202 800
rect 96434 0 96490 800
rect 97722 0 97778 800
rect 99010 0 99066 800
rect 100390 0 100446 800
rect 101678 0 101734 800
rect 102966 0 103022 800
rect 104254 0 104310 800
rect 105634 0 105690 800
rect 106922 0 106978 800
rect 108210 0 108266 800
rect 109498 0 109554 800
rect 110878 0 110934 800
rect 112166 0 112222 800
rect 113454 0 113510 800
rect 114834 0 114890 800
rect 116122 0 116178 800
rect 117410 0 117466 800
rect 118698 0 118754 800
rect 120078 0 120134 800
rect 121366 0 121422 800
rect 122654 0 122710 800
rect 123942 0 123998 800
rect 125322 0 125378 800
rect 126610 0 126666 800
rect 127898 0 127954 800
rect 129186 0 129242 800
rect 130566 0 130622 800
rect 131854 0 131910 800
rect 133142 0 133198 800
rect 134522 0 134578 800
rect 135810 0 135866 800
rect 137098 0 137154 800
rect 138386 0 138442 800
rect 139766 0 139822 800
rect 141054 0 141110 800
rect 142342 0 142398 800
rect 143630 0 143686 800
rect 145010 0 145066 800
rect 146298 0 146354 800
rect 147586 0 147642 800
rect 148874 0 148930 800
rect 150254 0 150310 800
rect 151542 0 151598 800
rect 152830 0 152886 800
rect 154118 0 154174 800
rect 155498 0 155554 800
rect 156786 0 156842 800
rect 158074 0 158130 800
rect 159454 0 159510 800
rect 160742 0 160798 800
rect 162030 0 162086 800
rect 163318 0 163374 800
rect 164698 0 164754 800
rect 165986 0 166042 800
rect 167274 0 167330 800
rect 168562 0 168618 800
rect 169942 0 169998 800
rect 171230 0 171286 800
rect 172518 0 172574 800
rect 173806 0 173862 800
rect 175186 0 175242 800
rect 176474 0 176530 800
rect 177762 0 177818 800
rect 179142 0 179198 800
rect 180430 0 180486 800
rect 181718 0 181774 800
rect 183006 0 183062 800
rect 184386 0 184442 800
rect 185674 0 185730 800
rect 186962 0 187018 800
rect 188250 0 188306 800
rect 189630 0 189686 800
rect 190918 0 190974 800
rect 192206 0 192262 800
rect 193494 0 193550 800
rect 194874 0 194930 800
rect 196162 0 196218 800
rect 197450 0 197506 800
<< obsm2 >>
rect 682 199448 1710 199594
rect 1878 199448 2998 199594
rect 3166 199448 4286 199594
rect 4454 199448 5574 199594
rect 5742 199448 6862 199594
rect 7030 199448 8150 199594
rect 8318 199448 9438 199594
rect 9606 199448 10726 199594
rect 10894 199448 12014 199594
rect 12182 199448 13210 199594
rect 13378 199448 14498 199594
rect 14666 199448 15786 199594
rect 15954 199448 17074 199594
rect 17242 199448 18362 199594
rect 18530 199448 19650 199594
rect 19818 199448 20938 199594
rect 21106 199448 22226 199594
rect 22394 199448 23514 199594
rect 23682 199448 24802 199594
rect 24970 199448 25998 199594
rect 26166 199448 27286 199594
rect 27454 199448 28574 199594
rect 28742 199448 29862 199594
rect 30030 199448 31150 199594
rect 31318 199448 32438 199594
rect 32606 199448 33726 199594
rect 33894 199448 35014 199594
rect 35182 199448 36302 199594
rect 36470 199448 37590 199594
rect 37758 199448 38786 199594
rect 38954 199448 40074 199594
rect 40242 199448 41362 199594
rect 41530 199448 42650 199594
rect 42818 199448 43938 199594
rect 44106 199448 45226 199594
rect 45394 199448 46514 199594
rect 46682 199448 47802 199594
rect 47970 199448 49090 199594
rect 49258 199448 50286 199594
rect 50454 199448 51574 199594
rect 51742 199448 52862 199594
rect 53030 199448 54150 199594
rect 54318 199448 55438 199594
rect 55606 199448 56726 199594
rect 56894 199448 58014 199594
rect 58182 199448 59302 199594
rect 59470 199448 60590 199594
rect 60758 199448 61878 199594
rect 62046 199448 63074 199594
rect 63242 199448 64362 199594
rect 64530 199448 65650 199594
rect 65818 199448 66938 199594
rect 67106 199448 68226 199594
rect 68394 199448 69514 199594
rect 69682 199448 70802 199594
rect 70970 199448 72090 199594
rect 72258 199448 73378 199594
rect 73546 199448 74666 199594
rect 74834 199448 75862 199594
rect 76030 199448 77150 199594
rect 77318 199448 78438 199594
rect 78606 199448 79726 199594
rect 79894 199448 81014 199594
rect 81182 199448 82302 199594
rect 82470 199448 83590 199594
rect 83758 199448 84878 199594
rect 85046 199448 86166 199594
rect 86334 199448 87362 199594
rect 87530 199448 88650 199594
rect 88818 199448 89938 199594
rect 90106 199448 91226 199594
rect 91394 199448 92514 199594
rect 92682 199448 93802 199594
rect 93970 199448 95090 199594
rect 95258 199448 96378 199594
rect 96546 199448 97666 199594
rect 97834 199448 98954 199594
rect 99122 199448 100150 199594
rect 100318 199448 101438 199594
rect 101606 199448 102726 199594
rect 102894 199448 104014 199594
rect 104182 199448 105302 199594
rect 105470 199448 106590 199594
rect 106758 199448 107878 199594
rect 108046 199448 109166 199594
rect 109334 199448 110454 199594
rect 110622 199448 111742 199594
rect 111910 199448 112938 199594
rect 113106 199448 114226 199594
rect 114394 199448 115514 199594
rect 115682 199448 116802 199594
rect 116970 199448 118090 199594
rect 118258 199448 119378 199594
rect 119546 199448 120666 199594
rect 120834 199448 121954 199594
rect 122122 199448 123242 199594
rect 123410 199448 124438 199594
rect 124606 199448 125726 199594
rect 125894 199448 127014 199594
rect 127182 199448 128302 199594
rect 128470 199448 129590 199594
rect 129758 199448 130878 199594
rect 131046 199448 132166 199594
rect 132334 199448 133454 199594
rect 133622 199448 134742 199594
rect 134910 199448 136030 199594
rect 136198 199448 137226 199594
rect 137394 199448 138514 199594
rect 138682 199448 139802 199594
rect 139970 199448 141090 199594
rect 141258 199448 142378 199594
rect 142546 199448 143666 199594
rect 143834 199448 144954 199594
rect 145122 199448 146242 199594
rect 146410 199448 147530 199594
rect 147698 199448 148818 199594
rect 148986 199448 150014 199594
rect 150182 199448 151302 199594
rect 151470 199448 152590 199594
rect 152758 199448 153878 199594
rect 154046 199448 155166 199594
rect 155334 199448 156454 199594
rect 156622 199448 157742 199594
rect 157910 199448 159030 199594
rect 159198 199448 160318 199594
rect 160486 199448 161514 199594
rect 161682 199448 162802 199594
rect 162970 199448 164090 199594
rect 164258 199448 165378 199594
rect 165546 199448 166666 199594
rect 166834 199448 167954 199594
rect 168122 199448 169242 199594
rect 169410 199448 170530 199594
rect 170698 199448 171818 199594
rect 171986 199448 173106 199594
rect 173274 199448 174302 199594
rect 174470 199448 175590 199594
rect 175758 199448 176878 199594
rect 177046 199448 178166 199594
rect 178334 199448 179454 199594
rect 179622 199448 180742 199594
rect 180910 199448 182030 199594
rect 182198 199448 183318 199594
rect 183486 199448 184606 199594
rect 184774 199448 185894 199594
rect 186062 199448 187090 199594
rect 187258 199448 188378 199594
rect 188546 199448 189666 199594
rect 189834 199448 190954 199594
rect 191122 199448 192242 199594
rect 192410 199448 193530 199594
rect 193698 199448 194818 199594
rect 194986 199448 196106 199594
rect 196274 199448 197394 199594
rect 676 856 197504 199448
rect 774 31 1894 856
rect 2062 31 3182 856
rect 3350 31 4470 856
rect 4638 31 5850 856
rect 6018 31 7138 856
rect 7306 31 8426 856
rect 8594 31 9714 856
rect 9882 31 11094 856
rect 11262 31 12382 856
rect 12550 31 13670 856
rect 13838 31 14958 856
rect 15126 31 16338 856
rect 16506 31 17626 856
rect 17794 31 18914 856
rect 19082 31 20202 856
rect 20370 31 21582 856
rect 21750 31 22870 856
rect 23038 31 24158 856
rect 24326 31 25538 856
rect 25706 31 26826 856
rect 26994 31 28114 856
rect 28282 31 29402 856
rect 29570 31 30782 856
rect 30950 31 32070 856
rect 32238 31 33358 856
rect 33526 31 34646 856
rect 34814 31 36026 856
rect 36194 31 37314 856
rect 37482 31 38602 856
rect 38770 31 39890 856
rect 40058 31 41270 856
rect 41438 31 42558 856
rect 42726 31 43846 856
rect 44014 31 45226 856
rect 45394 31 46514 856
rect 46682 31 47802 856
rect 47970 31 49090 856
rect 49258 31 50470 856
rect 50638 31 51758 856
rect 51926 31 53046 856
rect 53214 31 54334 856
rect 54502 31 55714 856
rect 55882 31 57002 856
rect 57170 31 58290 856
rect 58458 31 59578 856
rect 59746 31 60958 856
rect 61126 31 62246 856
rect 62414 31 63534 856
rect 63702 31 64822 856
rect 64990 31 66202 856
rect 66370 31 67490 856
rect 67658 31 68778 856
rect 68946 31 70158 856
rect 70326 31 71446 856
rect 71614 31 72734 856
rect 72902 31 74022 856
rect 74190 31 75402 856
rect 75570 31 76690 856
rect 76858 31 77978 856
rect 78146 31 79266 856
rect 79434 31 80646 856
rect 80814 31 81934 856
rect 82102 31 83222 856
rect 83390 31 84510 856
rect 84678 31 85890 856
rect 86058 31 87178 856
rect 87346 31 88466 856
rect 88634 31 89846 856
rect 90014 31 91134 856
rect 91302 31 92422 856
rect 92590 31 93710 856
rect 93878 31 95090 856
rect 95258 31 96378 856
rect 96546 31 97666 856
rect 97834 31 98954 856
rect 99122 31 100334 856
rect 100502 31 101622 856
rect 101790 31 102910 856
rect 103078 31 104198 856
rect 104366 31 105578 856
rect 105746 31 106866 856
rect 107034 31 108154 856
rect 108322 31 109442 856
rect 109610 31 110822 856
rect 110990 31 112110 856
rect 112278 31 113398 856
rect 113566 31 114778 856
rect 114946 31 116066 856
rect 116234 31 117354 856
rect 117522 31 118642 856
rect 118810 31 120022 856
rect 120190 31 121310 856
rect 121478 31 122598 856
rect 122766 31 123886 856
rect 124054 31 125266 856
rect 125434 31 126554 856
rect 126722 31 127842 856
rect 128010 31 129130 856
rect 129298 31 130510 856
rect 130678 31 131798 856
rect 131966 31 133086 856
rect 133254 31 134466 856
rect 134634 31 135754 856
rect 135922 31 137042 856
rect 137210 31 138330 856
rect 138498 31 139710 856
rect 139878 31 140998 856
rect 141166 31 142286 856
rect 142454 31 143574 856
rect 143742 31 144954 856
rect 145122 31 146242 856
rect 146410 31 147530 856
rect 147698 31 148818 856
rect 148986 31 150198 856
rect 150366 31 151486 856
rect 151654 31 152774 856
rect 152942 31 154062 856
rect 154230 31 155442 856
rect 155610 31 156730 856
rect 156898 31 158018 856
rect 158186 31 159398 856
rect 159566 31 160686 856
rect 160854 31 161974 856
rect 162142 31 163262 856
rect 163430 31 164642 856
rect 164810 31 165930 856
rect 166098 31 167218 856
rect 167386 31 168506 856
rect 168674 31 169886 856
rect 170054 31 171174 856
rect 171342 31 172462 856
rect 172630 31 173750 856
rect 173918 31 175130 856
rect 175298 31 176418 856
rect 176586 31 177706 856
rect 177874 31 179086 856
rect 179254 31 180374 856
rect 180542 31 181662 856
rect 181830 31 182950 856
rect 183118 31 184330 856
rect 184498 31 185618 856
rect 185786 31 186906 856
rect 187074 31 188194 856
rect 188362 31 189574 856
rect 189742 31 190862 856
rect 191030 31 192150 856
rect 192318 31 193438 856
rect 193606 31 194818 856
rect 194986 31 196106 856
rect 196274 31 197394 856
<< metal3 >>
rect 197360 197752 198160 197872
rect 0 197480 800 197600
rect 197360 192720 198160 192840
rect 0 192040 800 192160
rect 197360 187688 198160 187808
rect 0 186600 800 186720
rect 197360 182656 198160 182776
rect 0 181160 800 181280
rect 197360 177624 198160 177744
rect 0 175720 800 175840
rect 197360 172728 198160 172848
rect 0 170416 800 170536
rect 197360 167696 198160 167816
rect 0 164976 800 165096
rect 197360 162664 198160 162784
rect 0 159536 800 159656
rect 197360 157632 198160 157752
rect 0 154096 800 154216
rect 197360 152600 198160 152720
rect 0 148656 800 148776
rect 197360 147568 198160 147688
rect 0 143352 800 143472
rect 197360 142672 198160 142792
rect 0 137912 800 138032
rect 197360 137640 198160 137760
rect 0 132472 800 132592
rect 197360 132608 198160 132728
rect 197360 127576 198160 127696
rect 0 127032 800 127152
rect 197360 122544 198160 122664
rect 0 121592 800 121712
rect 197360 117512 198160 117632
rect 0 116288 800 116408
rect 197360 112616 198160 112736
rect 0 110848 800 110968
rect 197360 107584 198160 107704
rect 0 105408 800 105528
rect 197360 102552 198160 102672
rect 0 99968 800 100088
rect 197360 97520 198160 97640
rect 0 94528 800 94648
rect 197360 92488 198160 92608
rect 0 89088 800 89208
rect 197360 87592 198160 87712
rect 0 83784 800 83904
rect 197360 82560 198160 82680
rect 0 78344 800 78464
rect 197360 77528 198160 77648
rect 0 72904 800 73024
rect 197360 72496 198160 72616
rect 0 67464 800 67584
rect 197360 67464 198160 67584
rect 197360 62432 198160 62552
rect 0 62024 800 62144
rect 197360 57536 198160 57656
rect 0 56720 800 56840
rect 197360 52504 198160 52624
rect 0 51280 800 51400
rect 197360 47472 198160 47592
rect 0 45840 800 45960
rect 197360 42440 198160 42560
rect 0 40400 800 40520
rect 197360 37408 198160 37528
rect 0 34960 800 35080
rect 197360 32376 198160 32496
rect 0 29656 800 29776
rect 197360 27480 198160 27600
rect 0 24216 800 24336
rect 197360 22448 198160 22568
rect 0 18776 800 18896
rect 197360 17416 198160 17536
rect 0 13336 800 13456
rect 197360 12384 198160 12504
rect 0 7896 800 8016
rect 197360 7352 198160 7472
rect 0 2592 800 2712
rect 197360 2456 198160 2576
<< obsm3 >>
rect 749 197952 197360 198253
rect 749 197680 197280 197952
rect 880 197672 197280 197680
rect 880 197400 197360 197672
rect 749 192920 197360 197400
rect 749 192640 197280 192920
rect 749 192240 197360 192640
rect 880 191960 197360 192240
rect 749 187888 197360 191960
rect 749 187608 197280 187888
rect 749 186800 197360 187608
rect 880 186520 197360 186800
rect 749 182856 197360 186520
rect 749 182576 197280 182856
rect 749 181360 197360 182576
rect 880 181080 197360 181360
rect 749 177824 197360 181080
rect 749 177544 197280 177824
rect 749 175920 197360 177544
rect 880 175640 197360 175920
rect 749 172928 197360 175640
rect 749 172648 197280 172928
rect 749 170616 197360 172648
rect 880 170336 197360 170616
rect 749 167896 197360 170336
rect 749 167616 197280 167896
rect 749 165176 197360 167616
rect 880 164896 197360 165176
rect 749 162864 197360 164896
rect 749 162584 197280 162864
rect 749 159736 197360 162584
rect 880 159456 197360 159736
rect 749 157832 197360 159456
rect 749 157552 197280 157832
rect 749 154296 197360 157552
rect 880 154016 197360 154296
rect 749 152800 197360 154016
rect 749 152520 197280 152800
rect 749 148856 197360 152520
rect 880 148576 197360 148856
rect 749 147768 197360 148576
rect 749 147488 197280 147768
rect 749 143552 197360 147488
rect 880 143272 197360 143552
rect 749 142872 197360 143272
rect 749 142592 197280 142872
rect 749 138112 197360 142592
rect 880 137840 197360 138112
rect 880 137832 197280 137840
rect 749 137560 197280 137832
rect 749 132808 197360 137560
rect 749 132672 197280 132808
rect 880 132528 197280 132672
rect 880 132392 197360 132528
rect 749 127776 197360 132392
rect 749 127496 197280 127776
rect 749 127232 197360 127496
rect 880 126952 197360 127232
rect 749 122744 197360 126952
rect 749 122464 197280 122744
rect 749 121792 197360 122464
rect 880 121512 197360 121792
rect 749 117712 197360 121512
rect 749 117432 197280 117712
rect 749 116488 197360 117432
rect 880 116208 197360 116488
rect 749 112816 197360 116208
rect 749 112536 197280 112816
rect 749 111048 197360 112536
rect 880 110768 197360 111048
rect 749 107784 197360 110768
rect 749 107504 197280 107784
rect 749 105608 197360 107504
rect 880 105328 197360 105608
rect 749 102752 197360 105328
rect 749 102472 197280 102752
rect 749 100168 197360 102472
rect 880 99888 197360 100168
rect 749 97720 197360 99888
rect 749 97440 197280 97720
rect 749 94728 197360 97440
rect 880 94448 197360 94728
rect 749 92688 197360 94448
rect 749 92408 197280 92688
rect 749 89288 197360 92408
rect 880 89008 197360 89288
rect 749 87792 197360 89008
rect 749 87512 197280 87792
rect 749 83984 197360 87512
rect 880 83704 197360 83984
rect 749 82760 197360 83704
rect 749 82480 197280 82760
rect 749 78544 197360 82480
rect 880 78264 197360 78544
rect 749 77728 197360 78264
rect 749 77448 197280 77728
rect 749 73104 197360 77448
rect 880 72824 197360 73104
rect 749 72696 197360 72824
rect 749 72416 197280 72696
rect 749 67664 197360 72416
rect 880 67384 197280 67664
rect 749 62632 197360 67384
rect 749 62352 197280 62632
rect 749 62224 197360 62352
rect 880 61944 197360 62224
rect 749 57736 197360 61944
rect 749 57456 197280 57736
rect 749 56920 197360 57456
rect 880 56640 197360 56920
rect 749 52704 197360 56640
rect 749 52424 197280 52704
rect 749 51480 197360 52424
rect 880 51200 197360 51480
rect 749 47672 197360 51200
rect 749 47392 197280 47672
rect 749 46040 197360 47392
rect 880 45760 197360 46040
rect 749 42640 197360 45760
rect 749 42360 197280 42640
rect 749 40600 197360 42360
rect 880 40320 197360 40600
rect 749 37608 197360 40320
rect 749 37328 197280 37608
rect 749 35160 197360 37328
rect 880 34880 197360 35160
rect 749 32576 197360 34880
rect 749 32296 197280 32576
rect 749 29856 197360 32296
rect 880 29576 197360 29856
rect 749 27680 197360 29576
rect 749 27400 197280 27680
rect 749 24416 197360 27400
rect 880 24136 197360 24416
rect 749 22648 197360 24136
rect 749 22368 197280 22648
rect 749 18976 197360 22368
rect 880 18696 197360 18976
rect 749 17616 197360 18696
rect 749 17336 197280 17616
rect 749 13536 197360 17336
rect 880 13256 197360 13536
rect 749 12584 197360 13256
rect 749 12304 197280 12584
rect 749 8096 197360 12304
rect 880 7816 197360 8096
rect 749 7552 197360 7816
rect 749 7272 197280 7552
rect 749 2792 197360 7272
rect 880 2656 197360 2792
rect 880 2512 197280 2656
rect 749 2376 197280 2512
rect 749 35 197360 2376
<< metal4 >>
rect 4208 2128 4528 198064
rect 19568 2128 19888 198064
rect 34928 2128 35248 198064
rect 50288 2128 50608 198064
rect 65648 2128 65968 198064
rect 81008 2128 81328 198064
rect 96368 2128 96688 198064
rect 111728 2128 112048 198064
rect 127088 2128 127408 198064
rect 142448 2128 142768 198064
rect 157808 2128 158128 198064
rect 173168 2128 173488 198064
rect 188528 2128 188848 198064
<< obsm4 >>
rect 20115 198144 191117 198253
rect 20115 2619 34848 198144
rect 35328 2619 50208 198144
rect 50688 2619 65568 198144
rect 66048 2619 80928 198144
rect 81408 2619 96288 198144
rect 96768 2619 111648 198144
rect 112128 2619 127008 198144
rect 127488 2619 142368 198144
rect 142848 2619 157728 198144
rect 158208 2619 173088 198144
rect 173568 2619 188448 198144
rect 188928 2619 191117 198144
<< labels >>
rlabel metal2 s 143630 0 143686 800 6 clk_i
port 1 nsew signal input
rlabel metal3 s 197360 2456 198160 2576 6 i_dout0[0]
port 2 nsew signal input
rlabel metal2 s 168010 199504 168066 200304 6 i_dout0[10]
port 3 nsew signal input
rlabel metal2 s 170586 199504 170642 200304 6 i_dout0[11]
port 4 nsew signal input
rlabel metal3 s 0 105408 800 105528 6 i_dout0[12]
port 5 nsew signal input
rlabel metal3 s 197360 107584 198160 107704 6 i_dout0[13]
port 6 nsew signal input
rlabel metal2 s 169942 0 169998 800 6 i_dout0[14]
port 7 nsew signal input
rlabel metal3 s 0 121592 800 121712 6 i_dout0[15]
port 8 nsew signal input
rlabel metal3 s 197360 127576 198160 127696 6 i_dout0[16]
port 9 nsew signal input
rlabel metal2 s 175186 0 175242 800 6 i_dout0[17]
port 10 nsew signal input
rlabel metal3 s 0 143352 800 143472 6 i_dout0[18]
port 11 nsew signal input
rlabel metal2 s 177762 0 177818 800 6 i_dout0[19]
port 12 nsew signal input
rlabel metal2 s 147586 0 147642 800 6 i_dout0[1]
port 13 nsew signal input
rlabel metal2 s 180430 0 180486 800 6 i_dout0[20]
port 14 nsew signal input
rlabel metal2 s 182086 199504 182142 200304 6 i_dout0[21]
port 15 nsew signal input
rlabel metal3 s 0 170416 800 170536 6 i_dout0[22]
port 16 nsew signal input
rlabel metal3 s 0 175720 800 175840 6 i_dout0[23]
port 17 nsew signal input
rlabel metal2 s 184662 199504 184718 200304 6 i_dout0[24]
port 18 nsew signal input
rlabel metal2 s 187146 199504 187202 200304 6 i_dout0[25]
port 19 nsew signal input
rlabel metal3 s 197360 177624 198160 177744 6 i_dout0[26]
port 20 nsew signal input
rlabel metal3 s 197360 187688 198160 187808 6 i_dout0[27]
port 21 nsew signal input
rlabel metal2 s 190918 0 190974 800 6 i_dout0[28]
port 22 nsew signal input
rlabel metal3 s 197360 192720 198160 192840 6 i_dout0[29]
port 23 nsew signal input
rlabel metal2 s 148874 0 148930 800 6 i_dout0[2]
port 24 nsew signal input
rlabel metal2 s 193494 0 193550 800 6 i_dout0[30]
port 25 nsew signal input
rlabel metal2 s 196162 0 196218 800 6 i_dout0[31]
port 26 nsew signal input
rlabel metal3 s 0 45840 800 45960 6 i_dout0[3]
port 27 nsew signal input
rlabel metal2 s 151542 0 151598 800 6 i_dout0[4]
port 28 nsew signal input
rlabel metal2 s 161570 199504 161626 200304 6 i_dout0[5]
port 29 nsew signal input
rlabel metal3 s 0 78344 800 78464 6 i_dout0[6]
port 30 nsew signal input
rlabel metal3 s 197360 77528 198160 77648 6 i_dout0[7]
port 31 nsew signal input
rlabel metal2 s 160742 0 160798 800 6 i_dout0[8]
port 32 nsew signal input
rlabel metal2 s 166722 199504 166778 200304 6 i_dout0[9]
port 33 nsew signal input
rlabel metal3 s 0 13336 800 13456 6 i_dout0_1[0]
port 34 nsew signal input
rlabel metal3 s 0 94528 800 94648 6 i_dout0_1[10]
port 35 nsew signal input
rlabel metal2 s 165986 0 166042 800 6 i_dout0_1[11]
port 36 nsew signal input
rlabel metal2 s 173162 199504 173218 200304 6 i_dout0_1[12]
port 37 nsew signal input
rlabel metal2 s 175646 199504 175702 200304 6 i_dout0_1[13]
port 38 nsew signal input
rlabel metal3 s 197360 117512 198160 117632 6 i_dout0_1[14]
port 39 nsew signal input
rlabel metal2 s 171230 0 171286 800 6 i_dout0_1[15]
port 40 nsew signal input
rlabel metal2 s 172518 0 172574 800 6 i_dout0_1[16]
port 41 nsew signal input
rlabel metal3 s 197360 132608 198160 132728 6 i_dout0_1[17]
port 42 nsew signal input
rlabel metal3 s 0 137912 800 138032 6 i_dout0_1[18]
port 43 nsew signal input
rlabel metal3 s 197360 142672 198160 142792 6 i_dout0_1[19]
port 44 nsew signal input
rlabel metal3 s 0 34960 800 35080 6 i_dout0_1[1]
port 45 nsew signal input
rlabel metal3 s 197360 147568 198160 147688 6 i_dout0_1[20]
port 46 nsew signal input
rlabel metal2 s 181718 0 181774 800 6 i_dout0_1[21]
port 47 nsew signal input
rlabel metal2 s 183006 0 183062 800 6 i_dout0_1[22]
port 48 nsew signal input
rlabel metal2 s 184386 0 184442 800 6 i_dout0_1[23]
port 49 nsew signal input
rlabel metal3 s 197360 162664 198160 162784 6 i_dout0_1[24]
port 50 nsew signal input
rlabel metal2 s 185950 199504 186006 200304 6 i_dout0_1[25]
port 51 nsew signal input
rlabel metal3 s 197360 172728 198160 172848 6 i_dout0_1[26]
port 52 nsew signal input
rlabel metal2 s 188250 0 188306 800 6 i_dout0_1[27]
port 53 nsew signal input
rlabel metal2 s 191010 199504 191066 200304 6 i_dout0_1[28]
port 54 nsew signal input
rlabel metal2 s 192206 0 192262 800 6 i_dout0_1[29]
port 55 nsew signal input
rlabel metal2 s 153934 199504 153990 200304 6 i_dout0_1[2]
port 56 nsew signal input
rlabel metal2 s 194874 199504 194930 200304 6 i_dout0_1[30]
port 57 nsew signal input
rlabel metal2 s 196162 199504 196218 200304 6 i_dout0_1[31]
port 58 nsew signal input
rlabel metal2 s 157798 199504 157854 200304 6 i_dout0_1[3]
port 59 nsew signal input
rlabel metal3 s 197360 52504 198160 52624 6 i_dout0_1[4]
port 60 nsew signal input
rlabel metal3 s 0 67464 800 67584 6 i_dout0_1[5]
port 61 nsew signal input
rlabel metal2 s 156786 0 156842 800 6 i_dout0_1[6]
port 62 nsew signal input
rlabel metal2 s 165434 199504 165490 200304 6 i_dout0_1[7]
port 63 nsew signal input
rlabel metal2 s 159454 0 159510 800 6 i_dout0_1[8]
port 64 nsew signal input
rlabel metal3 s 197360 97520 198160 97640 6 i_dout0_1[9]
port 65 nsew signal input
rlabel metal2 s 570 199504 626 200304 6 io_in[0]
port 66 nsew signal input
rlabel metal2 s 38842 199504 38898 200304 6 io_in[10]
port 67 nsew signal input
rlabel metal2 s 42706 199504 42762 200304 6 io_in[11]
port 68 nsew signal input
rlabel metal2 s 46570 199504 46626 200304 6 io_in[12]
port 69 nsew signal input
rlabel metal2 s 50342 199504 50398 200304 6 io_in[13]
port 70 nsew signal input
rlabel metal2 s 54206 199504 54262 200304 6 io_in[14]
port 71 nsew signal input
rlabel metal2 s 58070 199504 58126 200304 6 io_in[15]
port 72 nsew signal input
rlabel metal2 s 61934 199504 61990 200304 6 io_in[16]
port 73 nsew signal input
rlabel metal2 s 65706 199504 65762 200304 6 io_in[17]
port 74 nsew signal input
rlabel metal2 s 69570 199504 69626 200304 6 io_in[18]
port 75 nsew signal input
rlabel metal2 s 73434 199504 73490 200304 6 io_in[19]
port 76 nsew signal input
rlabel metal2 s 4342 199504 4398 200304 6 io_in[1]
port 77 nsew signal input
rlabel metal2 s 77206 199504 77262 200304 6 io_in[20]
port 78 nsew signal input
rlabel metal2 s 81070 199504 81126 200304 6 io_in[21]
port 79 nsew signal input
rlabel metal2 s 84934 199504 84990 200304 6 io_in[22]
port 80 nsew signal input
rlabel metal2 s 88706 199504 88762 200304 6 io_in[23]
port 81 nsew signal input
rlabel metal2 s 92570 199504 92626 200304 6 io_in[24]
port 82 nsew signal input
rlabel metal2 s 96434 199504 96490 200304 6 io_in[25]
port 83 nsew signal input
rlabel metal2 s 100206 199504 100262 200304 6 io_in[26]
port 84 nsew signal input
rlabel metal2 s 104070 199504 104126 200304 6 io_in[27]
port 85 nsew signal input
rlabel metal2 s 107934 199504 107990 200304 6 io_in[28]
port 86 nsew signal input
rlabel metal2 s 111798 199504 111854 200304 6 io_in[29]
port 87 nsew signal input
rlabel metal2 s 8206 199504 8262 200304 6 io_in[2]
port 88 nsew signal input
rlabel metal2 s 115570 199504 115626 200304 6 io_in[30]
port 89 nsew signal input
rlabel metal2 s 119434 199504 119490 200304 6 io_in[31]
port 90 nsew signal input
rlabel metal2 s 123298 199504 123354 200304 6 io_in[32]
port 91 nsew signal input
rlabel metal2 s 127070 199504 127126 200304 6 io_in[33]
port 92 nsew signal input
rlabel metal2 s 130934 199504 130990 200304 6 io_in[34]
port 93 nsew signal input
rlabel metal2 s 134798 199504 134854 200304 6 io_in[35]
port 94 nsew signal input
rlabel metal2 s 138570 199504 138626 200304 6 io_in[36]
port 95 nsew signal input
rlabel metal2 s 142434 199504 142490 200304 6 io_in[37]
port 96 nsew signal input
rlabel metal2 s 12070 199504 12126 200304 6 io_in[3]
port 97 nsew signal input
rlabel metal2 s 15842 199504 15898 200304 6 io_in[4]
port 98 nsew signal input
rlabel metal2 s 19706 199504 19762 200304 6 io_in[5]
port 99 nsew signal input
rlabel metal2 s 23570 199504 23626 200304 6 io_in[6]
port 100 nsew signal input
rlabel metal2 s 27342 199504 27398 200304 6 io_in[7]
port 101 nsew signal input
rlabel metal2 s 31206 199504 31262 200304 6 io_in[8]
port 102 nsew signal input
rlabel metal2 s 35070 199504 35126 200304 6 io_in[9]
port 103 nsew signal input
rlabel metal2 s 1766 199504 1822 200304 6 io_oeb[0]
port 104 nsew signal output
rlabel metal2 s 40130 199504 40186 200304 6 io_oeb[10]
port 105 nsew signal output
rlabel metal2 s 43994 199504 44050 200304 6 io_oeb[11]
port 106 nsew signal output
rlabel metal2 s 47858 199504 47914 200304 6 io_oeb[12]
port 107 nsew signal output
rlabel metal2 s 51630 199504 51686 200304 6 io_oeb[13]
port 108 nsew signal output
rlabel metal2 s 55494 199504 55550 200304 6 io_oeb[14]
port 109 nsew signal output
rlabel metal2 s 59358 199504 59414 200304 6 io_oeb[15]
port 110 nsew signal output
rlabel metal2 s 63130 199504 63186 200304 6 io_oeb[16]
port 111 nsew signal output
rlabel metal2 s 66994 199504 67050 200304 6 io_oeb[17]
port 112 nsew signal output
rlabel metal2 s 70858 199504 70914 200304 6 io_oeb[18]
port 113 nsew signal output
rlabel metal2 s 74722 199504 74778 200304 6 io_oeb[19]
port 114 nsew signal output
rlabel metal2 s 5630 199504 5686 200304 6 io_oeb[1]
port 115 nsew signal output
rlabel metal2 s 78494 199504 78550 200304 6 io_oeb[20]
port 116 nsew signal output
rlabel metal2 s 82358 199504 82414 200304 6 io_oeb[21]
port 117 nsew signal output
rlabel metal2 s 86222 199504 86278 200304 6 io_oeb[22]
port 118 nsew signal output
rlabel metal2 s 89994 199504 90050 200304 6 io_oeb[23]
port 119 nsew signal output
rlabel metal2 s 93858 199504 93914 200304 6 io_oeb[24]
port 120 nsew signal output
rlabel metal2 s 97722 199504 97778 200304 6 io_oeb[25]
port 121 nsew signal output
rlabel metal2 s 101494 199504 101550 200304 6 io_oeb[26]
port 122 nsew signal output
rlabel metal2 s 105358 199504 105414 200304 6 io_oeb[27]
port 123 nsew signal output
rlabel metal2 s 109222 199504 109278 200304 6 io_oeb[28]
port 124 nsew signal output
rlabel metal2 s 112994 199504 113050 200304 6 io_oeb[29]
port 125 nsew signal output
rlabel metal2 s 9494 199504 9550 200304 6 io_oeb[2]
port 126 nsew signal output
rlabel metal2 s 116858 199504 116914 200304 6 io_oeb[30]
port 127 nsew signal output
rlabel metal2 s 120722 199504 120778 200304 6 io_oeb[31]
port 128 nsew signal output
rlabel metal2 s 124494 199504 124550 200304 6 io_oeb[32]
port 129 nsew signal output
rlabel metal2 s 128358 199504 128414 200304 6 io_oeb[33]
port 130 nsew signal output
rlabel metal2 s 132222 199504 132278 200304 6 io_oeb[34]
port 131 nsew signal output
rlabel metal2 s 136086 199504 136142 200304 6 io_oeb[35]
port 132 nsew signal output
rlabel metal2 s 139858 199504 139914 200304 6 io_oeb[36]
port 133 nsew signal output
rlabel metal2 s 143722 199504 143778 200304 6 io_oeb[37]
port 134 nsew signal output
rlabel metal2 s 13266 199504 13322 200304 6 io_oeb[3]
port 135 nsew signal output
rlabel metal2 s 17130 199504 17186 200304 6 io_oeb[4]
port 136 nsew signal output
rlabel metal2 s 20994 199504 21050 200304 6 io_oeb[5]
port 137 nsew signal output
rlabel metal2 s 24858 199504 24914 200304 6 io_oeb[6]
port 138 nsew signal output
rlabel metal2 s 28630 199504 28686 200304 6 io_oeb[7]
port 139 nsew signal output
rlabel metal2 s 32494 199504 32550 200304 6 io_oeb[8]
port 140 nsew signal output
rlabel metal2 s 36358 199504 36414 200304 6 io_oeb[9]
port 141 nsew signal output
rlabel metal2 s 3054 199504 3110 200304 6 io_out[0]
port 142 nsew signal output
rlabel metal2 s 41418 199504 41474 200304 6 io_out[10]
port 143 nsew signal output
rlabel metal2 s 45282 199504 45338 200304 6 io_out[11]
port 144 nsew signal output
rlabel metal2 s 49146 199504 49202 200304 6 io_out[12]
port 145 nsew signal output
rlabel metal2 s 52918 199504 52974 200304 6 io_out[13]
port 146 nsew signal output
rlabel metal2 s 56782 199504 56838 200304 6 io_out[14]
port 147 nsew signal output
rlabel metal2 s 60646 199504 60702 200304 6 io_out[15]
port 148 nsew signal output
rlabel metal2 s 64418 199504 64474 200304 6 io_out[16]
port 149 nsew signal output
rlabel metal2 s 68282 199504 68338 200304 6 io_out[17]
port 150 nsew signal output
rlabel metal2 s 72146 199504 72202 200304 6 io_out[18]
port 151 nsew signal output
rlabel metal2 s 75918 199504 75974 200304 6 io_out[19]
port 152 nsew signal output
rlabel metal2 s 6918 199504 6974 200304 6 io_out[1]
port 153 nsew signal output
rlabel metal2 s 79782 199504 79838 200304 6 io_out[20]
port 154 nsew signal output
rlabel metal2 s 83646 199504 83702 200304 6 io_out[21]
port 155 nsew signal output
rlabel metal2 s 87418 199504 87474 200304 6 io_out[22]
port 156 nsew signal output
rlabel metal2 s 91282 199504 91338 200304 6 io_out[23]
port 157 nsew signal output
rlabel metal2 s 95146 199504 95202 200304 6 io_out[24]
port 158 nsew signal output
rlabel metal2 s 99010 199504 99066 200304 6 io_out[25]
port 159 nsew signal output
rlabel metal2 s 102782 199504 102838 200304 6 io_out[26]
port 160 nsew signal output
rlabel metal2 s 106646 199504 106702 200304 6 io_out[27]
port 161 nsew signal output
rlabel metal2 s 110510 199504 110566 200304 6 io_out[28]
port 162 nsew signal output
rlabel metal2 s 114282 199504 114338 200304 6 io_out[29]
port 163 nsew signal output
rlabel metal2 s 10782 199504 10838 200304 6 io_out[2]
port 164 nsew signal output
rlabel metal2 s 118146 199504 118202 200304 6 io_out[30]
port 165 nsew signal output
rlabel metal2 s 122010 199504 122066 200304 6 io_out[31]
port 166 nsew signal output
rlabel metal2 s 125782 199504 125838 200304 6 io_out[32]
port 167 nsew signal output
rlabel metal2 s 129646 199504 129702 200304 6 io_out[33]
port 168 nsew signal output
rlabel metal2 s 133510 199504 133566 200304 6 io_out[34]
port 169 nsew signal output
rlabel metal2 s 137282 199504 137338 200304 6 io_out[35]
port 170 nsew signal output
rlabel metal2 s 141146 199504 141202 200304 6 io_out[36]
port 171 nsew signal output
rlabel metal2 s 145010 199504 145066 200304 6 io_out[37]
port 172 nsew signal output
rlabel metal2 s 14554 199504 14610 200304 6 io_out[3]
port 173 nsew signal output
rlabel metal2 s 18418 199504 18474 200304 6 io_out[4]
port 174 nsew signal output
rlabel metal2 s 22282 199504 22338 200304 6 io_out[5]
port 175 nsew signal output
rlabel metal2 s 26054 199504 26110 200304 6 io_out[6]
port 176 nsew signal output
rlabel metal2 s 29918 199504 29974 200304 6 io_out[7]
port 177 nsew signal output
rlabel metal2 s 33782 199504 33838 200304 6 io_out[8]
port 178 nsew signal output
rlabel metal2 s 37646 199504 37702 200304 6 io_out[9]
port 179 nsew signal output
rlabel metal2 s 139766 0 139822 800 6 irq[0]
port 180 nsew signal output
rlabel metal2 s 141054 0 141110 800 6 irq[1]
port 181 nsew signal output
rlabel metal2 s 142342 0 142398 800 6 irq[2]
port 182 nsew signal output
rlabel metal3 s 0 2592 800 2712 6 o_csb0
port 183 nsew signal output
rlabel metal2 s 145010 0 145066 800 6 o_csb0_1
port 184 nsew signal output
rlabel metal3 s 0 18776 800 18896 6 o_din0[0]
port 185 nsew signal output
rlabel metal3 s 0 99968 800 100088 6 o_din0[10]
port 186 nsew signal output
rlabel metal2 s 167274 0 167330 800 6 o_din0[11]
port 187 nsew signal output
rlabel metal2 s 174358 199504 174414 200304 6 o_din0[12]
port 188 nsew signal output
rlabel metal3 s 197360 112616 198160 112736 6 o_din0[13]
port 189 nsew signal output
rlabel metal3 s 197360 122544 198160 122664 6 o_din0[14]
port 190 nsew signal output
rlabel metal2 s 176934 199504 176990 200304 6 o_din0[15]
port 191 nsew signal output
rlabel metal2 s 178222 199504 178278 200304 6 o_din0[16]
port 192 nsew signal output
rlabel metal2 s 176474 0 176530 800 6 o_din0[17]
port 193 nsew signal output
rlabel metal3 s 197360 137640 198160 137760 6 o_din0[18]
port 194 nsew signal output
rlabel metal2 s 179510 199504 179566 200304 6 o_din0[19]
port 195 nsew signal output
rlabel metal3 s 197360 17416 198160 17536 6 o_din0[1]
port 196 nsew signal output
rlabel metal3 s 0 154096 800 154216 6 o_din0[20]
port 197 nsew signal output
rlabel metal3 s 0 164976 800 165096 6 o_din0[21]
port 198 nsew signal output
rlabel metal3 s 197360 152600 198160 152720 6 o_din0[22]
port 199 nsew signal output
rlabel metal3 s 0 181160 800 181280 6 o_din0[23]
port 200 nsew signal output
rlabel metal2 s 186962 0 187018 800 6 o_din0[24]
port 201 nsew signal output
rlabel metal3 s 0 186600 800 186720 6 o_din0[25]
port 202 nsew signal output
rlabel metal3 s 197360 182656 198160 182776 6 o_din0[26]
port 203 nsew signal output
rlabel metal2 s 189722 199504 189778 200304 6 o_din0[27]
port 204 nsew signal output
rlabel metal2 s 192298 199504 192354 200304 6 o_din0[28]
port 205 nsew signal output
rlabel metal3 s 0 197480 800 197600 6 o_din0[29]
port 206 nsew signal output
rlabel metal3 s 197360 32376 198160 32496 6 o_din0[2]
port 207 nsew signal output
rlabel metal2 s 194874 0 194930 800 6 o_din0[30]
port 208 nsew signal output
rlabel metal2 s 197450 0 197506 800 6 o_din0[31]
port 209 nsew signal output
rlabel metal3 s 197360 42440 198160 42560 6 o_din0[3]
port 210 nsew signal output
rlabel metal2 s 152830 0 152886 800 6 o_din0[4]
port 211 nsew signal output
rlabel metal3 s 197360 57536 198160 57656 6 o_din0[5]
port 212 nsew signal output
rlabel metal2 s 162858 199504 162914 200304 6 o_din0[6]
port 213 nsew signal output
rlabel metal3 s 197360 82560 198160 82680 6 o_din0[7]
port 214 nsew signal output
rlabel metal2 s 163318 0 163374 800 6 o_din0[8]
port 215 nsew signal output
rlabel metal2 s 164698 0 164754 800 6 o_din0[9]
port 216 nsew signal output
rlabel metal2 s 148874 199504 148930 200304 6 o_din0_1[0]
port 217 nsew signal output
rlabel metal2 s 169298 199504 169354 200304 6 o_din0_1[10]
port 218 nsew signal output
rlabel metal2 s 171874 199504 171930 200304 6 o_din0_1[11]
port 219 nsew signal output
rlabel metal2 s 168562 0 168618 800 6 o_din0_1[12]
port 220 nsew signal output
rlabel metal3 s 0 110848 800 110968 6 o_din0_1[13]
port 221 nsew signal output
rlabel metal3 s 0 116288 800 116408 6 o_din0_1[14]
port 222 nsew signal output
rlabel metal3 s 0 127032 800 127152 6 o_din0_1[15]
port 223 nsew signal output
rlabel metal2 s 173806 0 173862 800 6 o_din0_1[16]
port 224 nsew signal output
rlabel metal3 s 0 132472 800 132592 6 o_din0_1[17]
port 225 nsew signal output
rlabel metal3 s 0 148656 800 148776 6 o_din0_1[18]
port 226 nsew signal output
rlabel metal2 s 179142 0 179198 800 6 o_din0_1[19]
port 227 nsew signal output
rlabel metal3 s 197360 12384 198160 12504 6 o_din0_1[1]
port 228 nsew signal output
rlabel metal2 s 180798 199504 180854 200304 6 o_din0_1[20]
port 229 nsew signal output
rlabel metal3 s 0 159536 800 159656 6 o_din0_1[21]
port 230 nsew signal output
rlabel metal2 s 183374 199504 183430 200304 6 o_din0_1[22]
port 231 nsew signal output
rlabel metal3 s 197360 157632 198160 157752 6 o_din0_1[23]
port 232 nsew signal output
rlabel metal2 s 185674 0 185730 800 6 o_din0_1[24]
port 233 nsew signal output
rlabel metal3 s 197360 167696 198160 167816 6 o_din0_1[25]
port 234 nsew signal output
rlabel metal2 s 188434 199504 188490 200304 6 o_din0_1[26]
port 235 nsew signal output
rlabel metal2 s 189630 0 189686 800 6 o_din0_1[27]
port 236 nsew signal output
rlabel metal3 s 0 192040 800 192160 6 o_din0_1[28]
port 237 nsew signal output
rlabel metal2 s 193586 199504 193642 200304 6 o_din0_1[29]
port 238 nsew signal output
rlabel metal3 s 197360 27480 198160 27600 6 o_din0_1[2]
port 239 nsew signal output
rlabel metal3 s 197360 197752 198160 197872 6 o_din0_1[30]
port 240 nsew signal output
rlabel metal2 s 197450 199504 197506 200304 6 o_din0_1[31]
port 241 nsew signal output
rlabel metal3 s 0 51280 800 51400 6 o_din0_1[3]
port 242 nsew signal output
rlabel metal2 s 160374 199504 160430 200304 6 o_din0_1[4]
port 243 nsew signal output
rlabel metal3 s 0 72904 800 73024 6 o_din0_1[5]
port 244 nsew signal output
rlabel metal3 s 197360 67464 198160 67584 6 o_din0_1[6]
port 245 nsew signal output
rlabel metal3 s 0 83784 800 83904 6 o_din0_1[7]
port 246 nsew signal output
rlabel metal2 s 162030 0 162086 800 6 o_din0_1[8]
port 247 nsew signal output
rlabel metal3 s 197360 102552 198160 102672 6 o_din0_1[9]
port 248 nsew signal output
rlabel metal3 s 197360 7352 198160 7472 6 o_waddr0[0]
port 249 nsew signal output
rlabel metal2 s 151358 199504 151414 200304 6 o_waddr0[1]
port 250 nsew signal output
rlabel metal2 s 156510 199504 156566 200304 6 o_waddr0[2]
port 251 nsew signal output
rlabel metal2 s 159086 199504 159142 200304 6 o_waddr0[3]
port 252 nsew signal output
rlabel metal3 s 0 62024 800 62144 6 o_waddr0[4]
port 253 nsew signal output
rlabel metal2 s 155498 0 155554 800 6 o_waddr0[5]
port 254 nsew signal output
rlabel metal2 s 164146 199504 164202 200304 6 o_waddr0[6]
port 255 nsew signal output
rlabel metal3 s 0 89088 800 89208 6 o_waddr0[7]
port 256 nsew signal output
rlabel metal3 s 197360 92488 198160 92608 6 o_waddr0[8]
port 257 nsew signal output
rlabel metal3 s 0 24216 800 24336 6 o_waddr0_1[0]
port 258 nsew signal output
rlabel metal2 s 150070 199504 150126 200304 6 o_waddr0_1[1]
port 259 nsew signal output
rlabel metal2 s 155222 199504 155278 200304 6 o_waddr0_1[2]
port 260 nsew signal output
rlabel metal2 s 150254 0 150310 800 6 o_waddr0_1[3]
port 261 nsew signal output
rlabel metal2 s 154118 0 154174 800 6 o_waddr0_1[4]
port 262 nsew signal output
rlabel metal3 s 197360 62432 198160 62552 6 o_waddr0_1[5]
port 263 nsew signal output
rlabel metal3 s 197360 72496 198160 72616 6 o_waddr0_1[6]
port 264 nsew signal output
rlabel metal2 s 158074 0 158130 800 6 o_waddr0_1[7]
port 265 nsew signal output
rlabel metal3 s 197360 87592 198160 87712 6 o_waddr0_1[8]
port 266 nsew signal output
rlabel metal2 s 146298 199504 146354 200304 6 o_web0
port 267 nsew signal output
rlabel metal2 s 147586 199504 147642 200304 6 o_web0_1
port 268 nsew signal output
rlabel metal2 s 146298 0 146354 800 6 o_wmask0[0]
port 269 nsew signal output
rlabel metal2 s 152646 199504 152702 200304 6 o_wmask0[1]
port 270 nsew signal output
rlabel metal3 s 0 40400 800 40520 6 o_wmask0[2]
port 271 nsew signal output
rlabel metal3 s 0 56720 800 56840 6 o_wmask0[3]
port 272 nsew signal output
rlabel metal3 s 0 29656 800 29776 6 o_wmask0_1[0]
port 273 nsew signal output
rlabel metal3 s 197360 22448 198160 22568 6 o_wmask0_1[1]
port 274 nsew signal output
rlabel metal3 s 197360 37408 198160 37528 6 o_wmask0_1[2]
port 275 nsew signal output
rlabel metal3 s 197360 47472 198160 47592 6 o_wmask0_1[3]
port 276 nsew signal output
rlabel metal3 s 0 7896 800 8016 6 rst_i
port 277 nsew signal input
rlabel metal4 s 4208 2128 4528 198064 6 vccd1
port 278 nsew power input
rlabel metal4 s 34928 2128 35248 198064 6 vccd1
port 278 nsew power input
rlabel metal4 s 65648 2128 65968 198064 6 vccd1
port 278 nsew power input
rlabel metal4 s 96368 2128 96688 198064 6 vccd1
port 278 nsew power input
rlabel metal4 s 127088 2128 127408 198064 6 vccd1
port 278 nsew power input
rlabel metal4 s 157808 2128 158128 198064 6 vccd1
port 278 nsew power input
rlabel metal4 s 188528 2128 188848 198064 6 vccd1
port 278 nsew power input
rlabel metal4 s 19568 2128 19888 198064 6 vssd1
port 279 nsew ground input
rlabel metal4 s 50288 2128 50608 198064 6 vssd1
port 279 nsew ground input
rlabel metal4 s 81008 2128 81328 198064 6 vssd1
port 279 nsew ground input
rlabel metal4 s 111728 2128 112048 198064 6 vssd1
port 279 nsew ground input
rlabel metal4 s 142448 2128 142768 198064 6 vssd1
port 279 nsew ground input
rlabel metal4 s 173168 2128 173488 198064 6 vssd1
port 279 nsew ground input
rlabel metal2 s 662 0 718 800 6 wb_clk_i
port 280 nsew signal input
rlabel metal2 s 1950 0 2006 800 6 wb_rst_i
port 281 nsew signal input
rlabel metal2 s 3238 0 3294 800 6 wbs_ack_o
port 282 nsew signal output
rlabel metal2 s 8482 0 8538 800 6 wbs_adr_i[0]
port 283 nsew signal input
rlabel metal2 s 53102 0 53158 800 6 wbs_adr_i[10]
port 284 nsew signal input
rlabel metal2 s 57058 0 57114 800 6 wbs_adr_i[11]
port 285 nsew signal input
rlabel metal2 s 61014 0 61070 800 6 wbs_adr_i[12]
port 286 nsew signal input
rlabel metal2 s 64878 0 64934 800 6 wbs_adr_i[13]
port 287 nsew signal input
rlabel metal2 s 68834 0 68890 800 6 wbs_adr_i[14]
port 288 nsew signal input
rlabel metal2 s 72790 0 72846 800 6 wbs_adr_i[15]
port 289 nsew signal input
rlabel metal2 s 76746 0 76802 800 6 wbs_adr_i[16]
port 290 nsew signal input
rlabel metal2 s 80702 0 80758 800 6 wbs_adr_i[17]
port 291 nsew signal input
rlabel metal2 s 84566 0 84622 800 6 wbs_adr_i[18]
port 292 nsew signal input
rlabel metal2 s 88522 0 88578 800 6 wbs_adr_i[19]
port 293 nsew signal input
rlabel metal2 s 13726 0 13782 800 6 wbs_adr_i[1]
port 294 nsew signal input
rlabel metal2 s 92478 0 92534 800 6 wbs_adr_i[20]
port 295 nsew signal input
rlabel metal2 s 96434 0 96490 800 6 wbs_adr_i[21]
port 296 nsew signal input
rlabel metal2 s 100390 0 100446 800 6 wbs_adr_i[22]
port 297 nsew signal input
rlabel metal2 s 104254 0 104310 800 6 wbs_adr_i[23]
port 298 nsew signal input
rlabel metal2 s 108210 0 108266 800 6 wbs_adr_i[24]
port 299 nsew signal input
rlabel metal2 s 112166 0 112222 800 6 wbs_adr_i[25]
port 300 nsew signal input
rlabel metal2 s 116122 0 116178 800 6 wbs_adr_i[26]
port 301 nsew signal input
rlabel metal2 s 120078 0 120134 800 6 wbs_adr_i[27]
port 302 nsew signal input
rlabel metal2 s 123942 0 123998 800 6 wbs_adr_i[28]
port 303 nsew signal input
rlabel metal2 s 127898 0 127954 800 6 wbs_adr_i[29]
port 304 nsew signal input
rlabel metal2 s 18970 0 19026 800 6 wbs_adr_i[2]
port 305 nsew signal input
rlabel metal2 s 131854 0 131910 800 6 wbs_adr_i[30]
port 306 nsew signal input
rlabel metal2 s 135810 0 135866 800 6 wbs_adr_i[31]
port 307 nsew signal input
rlabel metal2 s 24214 0 24270 800 6 wbs_adr_i[3]
port 308 nsew signal input
rlabel metal2 s 29458 0 29514 800 6 wbs_adr_i[4]
port 309 nsew signal input
rlabel metal2 s 33414 0 33470 800 6 wbs_adr_i[5]
port 310 nsew signal input
rlabel metal2 s 37370 0 37426 800 6 wbs_adr_i[6]
port 311 nsew signal input
rlabel metal2 s 41326 0 41382 800 6 wbs_adr_i[7]
port 312 nsew signal input
rlabel metal2 s 45282 0 45338 800 6 wbs_adr_i[8]
port 313 nsew signal input
rlabel metal2 s 49146 0 49202 800 6 wbs_adr_i[9]
port 314 nsew signal input
rlabel metal2 s 4526 0 4582 800 6 wbs_cyc_i
port 315 nsew signal input
rlabel metal2 s 9770 0 9826 800 6 wbs_dat_i[0]
port 316 nsew signal input
rlabel metal2 s 54390 0 54446 800 6 wbs_dat_i[10]
port 317 nsew signal input
rlabel metal2 s 58346 0 58402 800 6 wbs_dat_i[11]
port 318 nsew signal input
rlabel metal2 s 62302 0 62358 800 6 wbs_dat_i[12]
port 319 nsew signal input
rlabel metal2 s 66258 0 66314 800 6 wbs_dat_i[13]
port 320 nsew signal input
rlabel metal2 s 70214 0 70270 800 6 wbs_dat_i[14]
port 321 nsew signal input
rlabel metal2 s 74078 0 74134 800 6 wbs_dat_i[15]
port 322 nsew signal input
rlabel metal2 s 78034 0 78090 800 6 wbs_dat_i[16]
port 323 nsew signal input
rlabel metal2 s 81990 0 82046 800 6 wbs_dat_i[17]
port 324 nsew signal input
rlabel metal2 s 85946 0 86002 800 6 wbs_dat_i[18]
port 325 nsew signal input
rlabel metal2 s 89902 0 89958 800 6 wbs_dat_i[19]
port 326 nsew signal input
rlabel metal2 s 15014 0 15070 800 6 wbs_dat_i[1]
port 327 nsew signal input
rlabel metal2 s 93766 0 93822 800 6 wbs_dat_i[20]
port 328 nsew signal input
rlabel metal2 s 97722 0 97778 800 6 wbs_dat_i[21]
port 329 nsew signal input
rlabel metal2 s 101678 0 101734 800 6 wbs_dat_i[22]
port 330 nsew signal input
rlabel metal2 s 105634 0 105690 800 6 wbs_dat_i[23]
port 331 nsew signal input
rlabel metal2 s 109498 0 109554 800 6 wbs_dat_i[24]
port 332 nsew signal input
rlabel metal2 s 113454 0 113510 800 6 wbs_dat_i[25]
port 333 nsew signal input
rlabel metal2 s 117410 0 117466 800 6 wbs_dat_i[26]
port 334 nsew signal input
rlabel metal2 s 121366 0 121422 800 6 wbs_dat_i[27]
port 335 nsew signal input
rlabel metal2 s 125322 0 125378 800 6 wbs_dat_i[28]
port 336 nsew signal input
rlabel metal2 s 129186 0 129242 800 6 wbs_dat_i[29]
port 337 nsew signal input
rlabel metal2 s 20258 0 20314 800 6 wbs_dat_i[2]
port 338 nsew signal input
rlabel metal2 s 133142 0 133198 800 6 wbs_dat_i[30]
port 339 nsew signal input
rlabel metal2 s 137098 0 137154 800 6 wbs_dat_i[31]
port 340 nsew signal input
rlabel metal2 s 25594 0 25650 800 6 wbs_dat_i[3]
port 341 nsew signal input
rlabel metal2 s 30838 0 30894 800 6 wbs_dat_i[4]
port 342 nsew signal input
rlabel metal2 s 34702 0 34758 800 6 wbs_dat_i[5]
port 343 nsew signal input
rlabel metal2 s 38658 0 38714 800 6 wbs_dat_i[6]
port 344 nsew signal input
rlabel metal2 s 42614 0 42670 800 6 wbs_dat_i[7]
port 345 nsew signal input
rlabel metal2 s 46570 0 46626 800 6 wbs_dat_i[8]
port 346 nsew signal input
rlabel metal2 s 50526 0 50582 800 6 wbs_dat_i[9]
port 347 nsew signal input
rlabel metal2 s 11150 0 11206 800 6 wbs_dat_o[0]
port 348 nsew signal output
rlabel metal2 s 55770 0 55826 800 6 wbs_dat_o[10]
port 349 nsew signal output
rlabel metal2 s 59634 0 59690 800 6 wbs_dat_o[11]
port 350 nsew signal output
rlabel metal2 s 63590 0 63646 800 6 wbs_dat_o[12]
port 351 nsew signal output
rlabel metal2 s 67546 0 67602 800 6 wbs_dat_o[13]
port 352 nsew signal output
rlabel metal2 s 71502 0 71558 800 6 wbs_dat_o[14]
port 353 nsew signal output
rlabel metal2 s 75458 0 75514 800 6 wbs_dat_o[15]
port 354 nsew signal output
rlabel metal2 s 79322 0 79378 800 6 wbs_dat_o[16]
port 355 nsew signal output
rlabel metal2 s 83278 0 83334 800 6 wbs_dat_o[17]
port 356 nsew signal output
rlabel metal2 s 87234 0 87290 800 6 wbs_dat_o[18]
port 357 nsew signal output
rlabel metal2 s 91190 0 91246 800 6 wbs_dat_o[19]
port 358 nsew signal output
rlabel metal2 s 16394 0 16450 800 6 wbs_dat_o[1]
port 359 nsew signal output
rlabel metal2 s 95146 0 95202 800 6 wbs_dat_o[20]
port 360 nsew signal output
rlabel metal2 s 99010 0 99066 800 6 wbs_dat_o[21]
port 361 nsew signal output
rlabel metal2 s 102966 0 103022 800 6 wbs_dat_o[22]
port 362 nsew signal output
rlabel metal2 s 106922 0 106978 800 6 wbs_dat_o[23]
port 363 nsew signal output
rlabel metal2 s 110878 0 110934 800 6 wbs_dat_o[24]
port 364 nsew signal output
rlabel metal2 s 114834 0 114890 800 6 wbs_dat_o[25]
port 365 nsew signal output
rlabel metal2 s 118698 0 118754 800 6 wbs_dat_o[26]
port 366 nsew signal output
rlabel metal2 s 122654 0 122710 800 6 wbs_dat_o[27]
port 367 nsew signal output
rlabel metal2 s 126610 0 126666 800 6 wbs_dat_o[28]
port 368 nsew signal output
rlabel metal2 s 130566 0 130622 800 6 wbs_dat_o[29]
port 369 nsew signal output
rlabel metal2 s 21638 0 21694 800 6 wbs_dat_o[2]
port 370 nsew signal output
rlabel metal2 s 134522 0 134578 800 6 wbs_dat_o[30]
port 371 nsew signal output
rlabel metal2 s 138386 0 138442 800 6 wbs_dat_o[31]
port 372 nsew signal output
rlabel metal2 s 26882 0 26938 800 6 wbs_dat_o[3]
port 373 nsew signal output
rlabel metal2 s 32126 0 32182 800 6 wbs_dat_o[4]
port 374 nsew signal output
rlabel metal2 s 36082 0 36138 800 6 wbs_dat_o[5]
port 375 nsew signal output
rlabel metal2 s 39946 0 40002 800 6 wbs_dat_o[6]
port 376 nsew signal output
rlabel metal2 s 43902 0 43958 800 6 wbs_dat_o[7]
port 377 nsew signal output
rlabel metal2 s 47858 0 47914 800 6 wbs_dat_o[8]
port 378 nsew signal output
rlabel metal2 s 51814 0 51870 800 6 wbs_dat_o[9]
port 379 nsew signal output
rlabel metal2 s 12438 0 12494 800 6 wbs_sel_i[0]
port 380 nsew signal input
rlabel metal2 s 17682 0 17738 800 6 wbs_sel_i[1]
port 381 nsew signal input
rlabel metal2 s 22926 0 22982 800 6 wbs_sel_i[2]
port 382 nsew signal input
rlabel metal2 s 28170 0 28226 800 6 wbs_sel_i[3]
port 383 nsew signal input
rlabel metal2 s 5906 0 5962 800 6 wbs_stb_i
port 384 nsew signal input
rlabel metal2 s 7194 0 7250 800 6 wbs_we_i
port 385 nsew signal input
<< properties >>
string LEFclass BLOCK
string FIXED_BBOX 0 0 198160 200304
string LEFview TRUE
string GDS_FILE /local/home/roman/projects/opencircuitdesign/shuttle5/caravel_mpw/openlane/user_proj/runs/user_proj/results/magic/user_proj.gds
string GDS_END 97904358
string GDS_START 1523166
<< end >>

