magic
tech sky130A
magscale 1 2
timestamp 1643866341
<< obsli1 >>
rect 1104 2159 197403 198033
<< obsm1 >>
rect 658 960 197694 198212
<< metal2 >>
rect 570 199469 626 200269
rect 1766 199469 1822 200269
rect 3054 199469 3110 200269
rect 4342 199469 4398 200269
rect 5630 199469 5686 200269
rect 6918 199469 6974 200269
rect 8206 199469 8262 200269
rect 9494 199469 9550 200269
rect 10782 199469 10838 200269
rect 12070 199469 12126 200269
rect 13266 199469 13322 200269
rect 14554 199469 14610 200269
rect 15842 199469 15898 200269
rect 17130 199469 17186 200269
rect 18418 199469 18474 200269
rect 19706 199469 19762 200269
rect 20994 199469 21050 200269
rect 22282 199469 22338 200269
rect 23570 199469 23626 200269
rect 24858 199469 24914 200269
rect 26054 199469 26110 200269
rect 27342 199469 27398 200269
rect 28630 199469 28686 200269
rect 29918 199469 29974 200269
rect 31206 199469 31262 200269
rect 32494 199469 32550 200269
rect 33782 199469 33838 200269
rect 35070 199469 35126 200269
rect 36358 199469 36414 200269
rect 37646 199469 37702 200269
rect 38842 199469 38898 200269
rect 40130 199469 40186 200269
rect 41418 199469 41474 200269
rect 42706 199469 42762 200269
rect 43994 199469 44050 200269
rect 45282 199469 45338 200269
rect 46570 199469 46626 200269
rect 47858 199469 47914 200269
rect 49146 199469 49202 200269
rect 50342 199469 50398 200269
rect 51630 199469 51686 200269
rect 52918 199469 52974 200269
rect 54206 199469 54262 200269
rect 55494 199469 55550 200269
rect 56782 199469 56838 200269
rect 58070 199469 58126 200269
rect 59358 199469 59414 200269
rect 60646 199469 60702 200269
rect 61934 199469 61990 200269
rect 63130 199469 63186 200269
rect 64418 199469 64474 200269
rect 65706 199469 65762 200269
rect 66994 199469 67050 200269
rect 68282 199469 68338 200269
rect 69570 199469 69626 200269
rect 70858 199469 70914 200269
rect 72146 199469 72202 200269
rect 73434 199469 73490 200269
rect 74722 199469 74778 200269
rect 75918 199469 75974 200269
rect 77206 199469 77262 200269
rect 78494 199469 78550 200269
rect 79782 199469 79838 200269
rect 81070 199469 81126 200269
rect 82358 199469 82414 200269
rect 83646 199469 83702 200269
rect 84934 199469 84990 200269
rect 86222 199469 86278 200269
rect 87418 199469 87474 200269
rect 88706 199469 88762 200269
rect 89994 199469 90050 200269
rect 91282 199469 91338 200269
rect 92570 199469 92626 200269
rect 93858 199469 93914 200269
rect 95146 199469 95202 200269
rect 96434 199469 96490 200269
rect 97722 199469 97778 200269
rect 99010 199469 99066 200269
rect 100206 199469 100262 200269
rect 101494 199469 101550 200269
rect 102782 199469 102838 200269
rect 104070 199469 104126 200269
rect 105358 199469 105414 200269
rect 106646 199469 106702 200269
rect 107934 199469 107990 200269
rect 109222 199469 109278 200269
rect 110510 199469 110566 200269
rect 111798 199469 111854 200269
rect 112994 199469 113050 200269
rect 114282 199469 114338 200269
rect 115570 199469 115626 200269
rect 116858 199469 116914 200269
rect 118146 199469 118202 200269
rect 119434 199469 119490 200269
rect 120722 199469 120778 200269
rect 122010 199469 122066 200269
rect 123298 199469 123354 200269
rect 124494 199469 124550 200269
rect 125782 199469 125838 200269
rect 127070 199469 127126 200269
rect 128358 199469 128414 200269
rect 129646 199469 129702 200269
rect 130934 199469 130990 200269
rect 132222 199469 132278 200269
rect 133510 199469 133566 200269
rect 134798 199469 134854 200269
rect 136086 199469 136142 200269
rect 137282 199469 137338 200269
rect 138570 199469 138626 200269
rect 139858 199469 139914 200269
rect 141146 199469 141202 200269
rect 142434 199469 142490 200269
rect 143722 199469 143778 200269
rect 145010 199469 145066 200269
rect 146298 199469 146354 200269
rect 147586 199469 147642 200269
rect 148874 199469 148930 200269
rect 150070 199469 150126 200269
rect 151358 199469 151414 200269
rect 152646 199469 152702 200269
rect 153934 199469 153990 200269
rect 155222 199469 155278 200269
rect 156510 199469 156566 200269
rect 157798 199469 157854 200269
rect 159086 199469 159142 200269
rect 160374 199469 160430 200269
rect 161570 199469 161626 200269
rect 162858 199469 162914 200269
rect 164146 199469 164202 200269
rect 165434 199469 165490 200269
rect 166722 199469 166778 200269
rect 168010 199469 168066 200269
rect 169298 199469 169354 200269
rect 170586 199469 170642 200269
rect 171874 199469 171930 200269
rect 173162 199469 173218 200269
rect 174358 199469 174414 200269
rect 175646 199469 175702 200269
rect 176934 199469 176990 200269
rect 178222 199469 178278 200269
rect 179510 199469 179566 200269
rect 180798 199469 180854 200269
rect 182086 199469 182142 200269
rect 183374 199469 183430 200269
rect 184662 199469 184718 200269
rect 185950 199469 186006 200269
rect 187146 199469 187202 200269
rect 188434 199469 188490 200269
rect 189722 199469 189778 200269
rect 191010 199469 191066 200269
rect 192298 199469 192354 200269
rect 193586 199469 193642 200269
rect 194874 199469 194930 200269
rect 196162 199469 196218 200269
rect 197450 199469 197506 200269
rect 662 0 718 800
rect 1950 0 2006 800
rect 3238 0 3294 800
rect 4526 0 4582 800
rect 5814 0 5870 800
rect 7102 0 7158 800
rect 8390 0 8446 800
rect 9678 0 9734 800
rect 10966 0 11022 800
rect 12254 0 12310 800
rect 13542 0 13598 800
rect 14830 0 14886 800
rect 16118 0 16174 800
rect 17498 0 17554 800
rect 18786 0 18842 800
rect 20074 0 20130 800
rect 21362 0 21418 800
rect 22650 0 22706 800
rect 23938 0 23994 800
rect 25226 0 25282 800
rect 26514 0 26570 800
rect 27802 0 27858 800
rect 29090 0 29146 800
rect 30378 0 30434 800
rect 31666 0 31722 800
rect 32954 0 33010 800
rect 34334 0 34390 800
rect 35622 0 35678 800
rect 36910 0 36966 800
rect 38198 0 38254 800
rect 39486 0 39542 800
rect 40774 0 40830 800
rect 42062 0 42118 800
rect 43350 0 43406 800
rect 44638 0 44694 800
rect 45926 0 45982 800
rect 47214 0 47270 800
rect 48502 0 48558 800
rect 49790 0 49846 800
rect 51170 0 51226 800
rect 52458 0 52514 800
rect 53746 0 53802 800
rect 55034 0 55090 800
rect 56322 0 56378 800
rect 57610 0 57666 800
rect 58898 0 58954 800
rect 60186 0 60242 800
rect 61474 0 61530 800
rect 62762 0 62818 800
rect 64050 0 64106 800
rect 65338 0 65394 800
rect 66718 0 66774 800
rect 68006 0 68062 800
rect 69294 0 69350 800
rect 70582 0 70638 800
rect 71870 0 71926 800
rect 73158 0 73214 800
rect 74446 0 74502 800
rect 75734 0 75790 800
rect 77022 0 77078 800
rect 78310 0 78366 800
rect 79598 0 79654 800
rect 80886 0 80942 800
rect 82174 0 82230 800
rect 83554 0 83610 800
rect 84842 0 84898 800
rect 86130 0 86186 800
rect 87418 0 87474 800
rect 88706 0 88762 800
rect 89994 0 90050 800
rect 91282 0 91338 800
rect 92570 0 92626 800
rect 93858 0 93914 800
rect 95146 0 95202 800
rect 96434 0 96490 800
rect 97722 0 97778 800
rect 99010 0 99066 800
rect 100390 0 100446 800
rect 101678 0 101734 800
rect 102966 0 103022 800
rect 104254 0 104310 800
rect 105542 0 105598 800
rect 106830 0 106886 800
rect 108118 0 108174 800
rect 109406 0 109462 800
rect 110694 0 110750 800
rect 111982 0 112038 800
rect 113270 0 113326 800
rect 114558 0 114614 800
rect 115846 0 115902 800
rect 117226 0 117282 800
rect 118514 0 118570 800
rect 119802 0 119858 800
rect 121090 0 121146 800
rect 122378 0 122434 800
rect 123666 0 123722 800
rect 124954 0 125010 800
rect 126242 0 126298 800
rect 127530 0 127586 800
rect 128818 0 128874 800
rect 130106 0 130162 800
rect 131394 0 131450 800
rect 132774 0 132830 800
rect 134062 0 134118 800
rect 135350 0 135406 800
rect 136638 0 136694 800
rect 137926 0 137982 800
rect 139214 0 139270 800
rect 140502 0 140558 800
rect 141790 0 141846 800
rect 143078 0 143134 800
rect 144366 0 144422 800
rect 145654 0 145710 800
rect 146942 0 146998 800
rect 148230 0 148286 800
rect 149610 0 149666 800
rect 150898 0 150954 800
rect 152186 0 152242 800
rect 153474 0 153530 800
rect 154762 0 154818 800
rect 156050 0 156106 800
rect 157338 0 157394 800
rect 158626 0 158682 800
rect 159914 0 159970 800
rect 161202 0 161258 800
rect 162490 0 162546 800
rect 163778 0 163834 800
rect 165066 0 165122 800
rect 166446 0 166502 800
rect 167734 0 167790 800
rect 169022 0 169078 800
rect 170310 0 170366 800
rect 171598 0 171654 800
rect 172886 0 172942 800
rect 174174 0 174230 800
rect 175462 0 175518 800
rect 176750 0 176806 800
rect 178038 0 178094 800
rect 179326 0 179382 800
rect 180614 0 180670 800
rect 181902 0 181958 800
rect 183282 0 183338 800
rect 184570 0 184626 800
rect 185858 0 185914 800
rect 187146 0 187202 800
rect 188434 0 188490 800
rect 189722 0 189778 800
rect 191010 0 191066 800
rect 192298 0 192354 800
rect 193586 0 193642 800
rect 194874 0 194930 800
rect 196162 0 196218 800
rect 197450 0 197506 800
<< obsm2 >>
rect 682 199413 1710 199469
rect 1878 199413 2998 199469
rect 3166 199413 4286 199469
rect 4454 199413 5574 199469
rect 5742 199413 6862 199469
rect 7030 199413 8150 199469
rect 8318 199413 9438 199469
rect 9606 199413 10726 199469
rect 10894 199413 12014 199469
rect 12182 199413 13210 199469
rect 13378 199413 14498 199469
rect 14666 199413 15786 199469
rect 15954 199413 17074 199469
rect 17242 199413 18362 199469
rect 18530 199413 19650 199469
rect 19818 199413 20938 199469
rect 21106 199413 22226 199469
rect 22394 199413 23514 199469
rect 23682 199413 24802 199469
rect 24970 199413 25998 199469
rect 26166 199413 27286 199469
rect 27454 199413 28574 199469
rect 28742 199413 29862 199469
rect 30030 199413 31150 199469
rect 31318 199413 32438 199469
rect 32606 199413 33726 199469
rect 33894 199413 35014 199469
rect 35182 199413 36302 199469
rect 36470 199413 37590 199469
rect 37758 199413 38786 199469
rect 38954 199413 40074 199469
rect 40242 199413 41362 199469
rect 41530 199413 42650 199469
rect 42818 199413 43938 199469
rect 44106 199413 45226 199469
rect 45394 199413 46514 199469
rect 46682 199413 47802 199469
rect 47970 199413 49090 199469
rect 49258 199413 50286 199469
rect 50454 199413 51574 199469
rect 51742 199413 52862 199469
rect 53030 199413 54150 199469
rect 54318 199413 55438 199469
rect 55606 199413 56726 199469
rect 56894 199413 58014 199469
rect 58182 199413 59302 199469
rect 59470 199413 60590 199469
rect 60758 199413 61878 199469
rect 62046 199413 63074 199469
rect 63242 199413 64362 199469
rect 64530 199413 65650 199469
rect 65818 199413 66938 199469
rect 67106 199413 68226 199469
rect 68394 199413 69514 199469
rect 69682 199413 70802 199469
rect 70970 199413 72090 199469
rect 72258 199413 73378 199469
rect 73546 199413 74666 199469
rect 74834 199413 75862 199469
rect 76030 199413 77150 199469
rect 77318 199413 78438 199469
rect 78606 199413 79726 199469
rect 79894 199413 81014 199469
rect 81182 199413 82302 199469
rect 82470 199413 83590 199469
rect 83758 199413 84878 199469
rect 85046 199413 86166 199469
rect 86334 199413 87362 199469
rect 87530 199413 88650 199469
rect 88818 199413 89938 199469
rect 90106 199413 91226 199469
rect 91394 199413 92514 199469
rect 92682 199413 93802 199469
rect 93970 199413 95090 199469
rect 95258 199413 96378 199469
rect 96546 199413 97666 199469
rect 97834 199413 98954 199469
rect 99122 199413 100150 199469
rect 100318 199413 101438 199469
rect 101606 199413 102726 199469
rect 102894 199413 104014 199469
rect 104182 199413 105302 199469
rect 105470 199413 106590 199469
rect 106758 199413 107878 199469
rect 108046 199413 109166 199469
rect 109334 199413 110454 199469
rect 110622 199413 111742 199469
rect 111910 199413 112938 199469
rect 113106 199413 114226 199469
rect 114394 199413 115514 199469
rect 115682 199413 116802 199469
rect 116970 199413 118090 199469
rect 118258 199413 119378 199469
rect 119546 199413 120666 199469
rect 120834 199413 121954 199469
rect 122122 199413 123242 199469
rect 123410 199413 124438 199469
rect 124606 199413 125726 199469
rect 125894 199413 127014 199469
rect 127182 199413 128302 199469
rect 128470 199413 129590 199469
rect 129758 199413 130878 199469
rect 131046 199413 132166 199469
rect 132334 199413 133454 199469
rect 133622 199413 134742 199469
rect 134910 199413 136030 199469
rect 136198 199413 137226 199469
rect 137394 199413 138514 199469
rect 138682 199413 139802 199469
rect 139970 199413 141090 199469
rect 141258 199413 142378 199469
rect 142546 199413 143666 199469
rect 143834 199413 144954 199469
rect 145122 199413 146242 199469
rect 146410 199413 147530 199469
rect 147698 199413 148818 199469
rect 148986 199413 150014 199469
rect 150182 199413 151302 199469
rect 151470 199413 152590 199469
rect 152758 199413 153878 199469
rect 154046 199413 155166 199469
rect 155334 199413 156454 199469
rect 156622 199413 157742 199469
rect 157910 199413 159030 199469
rect 159198 199413 160318 199469
rect 160486 199413 161514 199469
rect 161682 199413 162802 199469
rect 162970 199413 164090 199469
rect 164258 199413 165378 199469
rect 165546 199413 166666 199469
rect 166834 199413 167954 199469
rect 168122 199413 169242 199469
rect 169410 199413 170530 199469
rect 170698 199413 171818 199469
rect 171986 199413 173106 199469
rect 173274 199413 174302 199469
rect 174470 199413 175590 199469
rect 175758 199413 176878 199469
rect 177046 199413 178166 199469
rect 178334 199413 179454 199469
rect 179622 199413 180742 199469
rect 180910 199413 182030 199469
rect 182198 199413 183318 199469
rect 183486 199413 184606 199469
rect 184774 199413 185894 199469
rect 186062 199413 187090 199469
rect 187258 199413 188378 199469
rect 188546 199413 189666 199469
rect 189834 199413 190954 199469
rect 191122 199413 192242 199469
rect 192410 199413 193530 199469
rect 193698 199413 194818 199469
rect 194986 199413 196106 199469
rect 196274 199413 197394 199469
rect 197562 199413 197690 199469
rect 664 856 197690 199413
rect 774 734 1894 856
rect 2062 734 3182 856
rect 3350 734 4470 856
rect 4638 734 5758 856
rect 5926 734 7046 856
rect 7214 734 8334 856
rect 8502 734 9622 856
rect 9790 734 10910 856
rect 11078 734 12198 856
rect 12366 734 13486 856
rect 13654 734 14774 856
rect 14942 734 16062 856
rect 16230 734 17442 856
rect 17610 734 18730 856
rect 18898 734 20018 856
rect 20186 734 21306 856
rect 21474 734 22594 856
rect 22762 734 23882 856
rect 24050 734 25170 856
rect 25338 734 26458 856
rect 26626 734 27746 856
rect 27914 734 29034 856
rect 29202 734 30322 856
rect 30490 734 31610 856
rect 31778 734 32898 856
rect 33066 734 34278 856
rect 34446 734 35566 856
rect 35734 734 36854 856
rect 37022 734 38142 856
rect 38310 734 39430 856
rect 39598 734 40718 856
rect 40886 734 42006 856
rect 42174 734 43294 856
rect 43462 734 44582 856
rect 44750 734 45870 856
rect 46038 734 47158 856
rect 47326 734 48446 856
rect 48614 734 49734 856
rect 49902 734 51114 856
rect 51282 734 52402 856
rect 52570 734 53690 856
rect 53858 734 54978 856
rect 55146 734 56266 856
rect 56434 734 57554 856
rect 57722 734 58842 856
rect 59010 734 60130 856
rect 60298 734 61418 856
rect 61586 734 62706 856
rect 62874 734 63994 856
rect 64162 734 65282 856
rect 65450 734 66662 856
rect 66830 734 67950 856
rect 68118 734 69238 856
rect 69406 734 70526 856
rect 70694 734 71814 856
rect 71982 734 73102 856
rect 73270 734 74390 856
rect 74558 734 75678 856
rect 75846 734 76966 856
rect 77134 734 78254 856
rect 78422 734 79542 856
rect 79710 734 80830 856
rect 80998 734 82118 856
rect 82286 734 83498 856
rect 83666 734 84786 856
rect 84954 734 86074 856
rect 86242 734 87362 856
rect 87530 734 88650 856
rect 88818 734 89938 856
rect 90106 734 91226 856
rect 91394 734 92514 856
rect 92682 734 93802 856
rect 93970 734 95090 856
rect 95258 734 96378 856
rect 96546 734 97666 856
rect 97834 734 98954 856
rect 99122 734 100334 856
rect 100502 734 101622 856
rect 101790 734 102910 856
rect 103078 734 104198 856
rect 104366 734 105486 856
rect 105654 734 106774 856
rect 106942 734 108062 856
rect 108230 734 109350 856
rect 109518 734 110638 856
rect 110806 734 111926 856
rect 112094 734 113214 856
rect 113382 734 114502 856
rect 114670 734 115790 856
rect 115958 734 117170 856
rect 117338 734 118458 856
rect 118626 734 119746 856
rect 119914 734 121034 856
rect 121202 734 122322 856
rect 122490 734 123610 856
rect 123778 734 124898 856
rect 125066 734 126186 856
rect 126354 734 127474 856
rect 127642 734 128762 856
rect 128930 734 130050 856
rect 130218 734 131338 856
rect 131506 734 132718 856
rect 132886 734 134006 856
rect 134174 734 135294 856
rect 135462 734 136582 856
rect 136750 734 137870 856
rect 138038 734 139158 856
rect 139326 734 140446 856
rect 140614 734 141734 856
rect 141902 734 143022 856
rect 143190 734 144310 856
rect 144478 734 145598 856
rect 145766 734 146886 856
rect 147054 734 148174 856
rect 148342 734 149554 856
rect 149722 734 150842 856
rect 151010 734 152130 856
rect 152298 734 153418 856
rect 153586 734 154706 856
rect 154874 734 155994 856
rect 156162 734 157282 856
rect 157450 734 158570 856
rect 158738 734 159858 856
rect 160026 734 161146 856
rect 161314 734 162434 856
rect 162602 734 163722 856
rect 163890 734 165010 856
rect 165178 734 166390 856
rect 166558 734 167678 856
rect 167846 734 168966 856
rect 169134 734 170254 856
rect 170422 734 171542 856
rect 171710 734 172830 856
rect 172998 734 174118 856
rect 174286 734 175406 856
rect 175574 734 176694 856
rect 176862 734 177982 856
rect 178150 734 179270 856
rect 179438 734 180558 856
rect 180726 734 181846 856
rect 182014 734 183226 856
rect 183394 734 184514 856
rect 184682 734 185802 856
rect 185970 734 187090 856
rect 187258 734 188378 856
rect 188546 734 189666 856
rect 189834 734 190954 856
rect 191122 734 192242 856
rect 192410 734 193530 856
rect 193698 734 194818 856
rect 194986 734 196106 856
rect 196274 734 197394 856
rect 197562 734 197690 856
<< metal3 >>
rect 0 197888 800 198008
rect 197325 196936 198125 197056
rect 0 193400 800 193520
rect 197325 190408 198125 190528
rect 0 188776 800 188896
rect 0 184288 800 184408
rect 197325 184016 198125 184136
rect 0 179664 800 179784
rect 197325 177488 198125 177608
rect 0 175176 800 175296
rect 197325 171096 198125 171216
rect 0 170552 800 170672
rect 0 166064 800 166184
rect 197325 164568 198125 164688
rect 0 161440 800 161560
rect 197325 158176 198125 158296
rect 0 156952 800 157072
rect 0 152328 800 152448
rect 197325 151648 198125 151768
rect 0 147840 800 147960
rect 197325 145256 198125 145376
rect 0 143216 800 143336
rect 0 138728 800 138848
rect 197325 138728 198125 138848
rect 0 134104 800 134224
rect 197325 132336 198125 132456
rect 0 129616 800 129736
rect 197325 125808 198125 125928
rect 0 124992 800 125112
rect 0 120504 800 120624
rect 197325 119416 198125 119536
rect 0 115880 800 116000
rect 197325 112888 198125 113008
rect 0 111392 800 111512
rect 0 106768 800 106888
rect 197325 106496 198125 106616
rect 0 102280 800 102400
rect 197325 99968 198125 100088
rect 0 97792 800 97912
rect 197325 93576 198125 93696
rect 0 93168 800 93288
rect 0 88680 800 88800
rect 197325 87048 198125 87168
rect 0 84056 800 84176
rect 197325 80656 198125 80776
rect 0 79568 800 79688
rect 0 74944 800 75064
rect 197325 74128 198125 74248
rect 0 70456 800 70576
rect 197325 67736 198125 67856
rect 0 65832 800 65952
rect 0 61344 800 61464
rect 197325 61208 198125 61328
rect 0 56720 800 56840
rect 197325 54816 198125 54936
rect 0 52232 800 52352
rect 197325 48288 198125 48408
rect 0 47608 800 47728
rect 0 43120 800 43240
rect 197325 41896 198125 42016
rect 0 38496 800 38616
rect 197325 35368 198125 35488
rect 0 34008 800 34128
rect 0 29384 800 29504
rect 197325 28976 198125 29096
rect 0 24896 800 25016
rect 197325 22448 198125 22568
rect 0 20272 800 20392
rect 197325 16056 198125 16176
rect 0 15784 800 15904
rect 0 11160 800 11280
rect 197325 9528 198125 9648
rect 0 6672 800 6792
rect 197325 3136 198125 3256
rect 0 2184 800 2304
<< obsm3 >>
rect 800 198088 197695 198389
rect 880 197808 197695 198088
rect 800 197136 197695 197808
rect 800 196856 197245 197136
rect 800 193600 197695 196856
rect 880 193320 197695 193600
rect 800 190608 197695 193320
rect 800 190328 197245 190608
rect 800 188976 197695 190328
rect 880 188696 197695 188976
rect 800 184488 197695 188696
rect 880 184216 197695 184488
rect 880 184208 197245 184216
rect 800 183936 197245 184208
rect 800 179864 197695 183936
rect 880 179584 197695 179864
rect 800 177688 197695 179584
rect 800 177408 197245 177688
rect 800 175376 197695 177408
rect 880 175096 197695 175376
rect 800 171296 197695 175096
rect 800 171016 197245 171296
rect 800 170752 197695 171016
rect 880 170472 197695 170752
rect 800 166264 197695 170472
rect 880 165984 197695 166264
rect 800 164768 197695 165984
rect 800 164488 197245 164768
rect 800 161640 197695 164488
rect 880 161360 197695 161640
rect 800 158376 197695 161360
rect 800 158096 197245 158376
rect 800 157152 197695 158096
rect 880 156872 197695 157152
rect 800 152528 197695 156872
rect 880 152248 197695 152528
rect 800 151848 197695 152248
rect 800 151568 197245 151848
rect 800 148040 197695 151568
rect 880 147760 197695 148040
rect 800 145456 197695 147760
rect 800 145176 197245 145456
rect 800 143416 197695 145176
rect 880 143136 197695 143416
rect 800 138928 197695 143136
rect 880 138648 197245 138928
rect 800 134304 197695 138648
rect 880 134024 197695 134304
rect 800 132536 197695 134024
rect 800 132256 197245 132536
rect 800 129816 197695 132256
rect 880 129536 197695 129816
rect 800 126008 197695 129536
rect 800 125728 197245 126008
rect 800 125192 197695 125728
rect 880 124912 197695 125192
rect 800 120704 197695 124912
rect 880 120424 197695 120704
rect 800 119616 197695 120424
rect 800 119336 197245 119616
rect 800 116080 197695 119336
rect 880 115800 197695 116080
rect 800 113088 197695 115800
rect 800 112808 197245 113088
rect 800 111592 197695 112808
rect 880 111312 197695 111592
rect 800 106968 197695 111312
rect 880 106696 197695 106968
rect 880 106688 197245 106696
rect 800 106416 197245 106688
rect 800 102480 197695 106416
rect 880 102200 197695 102480
rect 800 100168 197695 102200
rect 800 99888 197245 100168
rect 800 97992 197695 99888
rect 880 97712 197695 97992
rect 800 93776 197695 97712
rect 800 93496 197245 93776
rect 800 93368 197695 93496
rect 880 93088 197695 93368
rect 800 88880 197695 93088
rect 880 88600 197695 88880
rect 800 87248 197695 88600
rect 800 86968 197245 87248
rect 800 84256 197695 86968
rect 880 83976 197695 84256
rect 800 80856 197695 83976
rect 800 80576 197245 80856
rect 800 79768 197695 80576
rect 880 79488 197695 79768
rect 800 75144 197695 79488
rect 880 74864 197695 75144
rect 800 74328 197695 74864
rect 800 74048 197245 74328
rect 800 70656 197695 74048
rect 880 70376 197695 70656
rect 800 67936 197695 70376
rect 800 67656 197245 67936
rect 800 66032 197695 67656
rect 880 65752 197695 66032
rect 800 61544 197695 65752
rect 880 61408 197695 61544
rect 880 61264 197245 61408
rect 800 61128 197245 61264
rect 800 56920 197695 61128
rect 880 56640 197695 56920
rect 800 55016 197695 56640
rect 800 54736 197245 55016
rect 800 52432 197695 54736
rect 880 52152 197695 52432
rect 800 48488 197695 52152
rect 800 48208 197245 48488
rect 800 47808 197695 48208
rect 880 47528 197695 47808
rect 800 43320 197695 47528
rect 880 43040 197695 43320
rect 800 42096 197695 43040
rect 800 41816 197245 42096
rect 800 38696 197695 41816
rect 880 38416 197695 38696
rect 800 35568 197695 38416
rect 800 35288 197245 35568
rect 800 34208 197695 35288
rect 880 33928 197695 34208
rect 800 29584 197695 33928
rect 880 29304 197695 29584
rect 800 29176 197695 29304
rect 800 28896 197245 29176
rect 800 25096 197695 28896
rect 880 24816 197695 25096
rect 800 22648 197695 24816
rect 800 22368 197245 22648
rect 800 20472 197695 22368
rect 880 20192 197695 20472
rect 800 16256 197695 20192
rect 800 15984 197245 16256
rect 880 15976 197245 15984
rect 880 15704 197695 15976
rect 800 11360 197695 15704
rect 880 11080 197695 11360
rect 800 9728 197695 11080
rect 800 9448 197245 9728
rect 800 6872 197695 9448
rect 880 6592 197695 6872
rect 800 3336 197695 6592
rect 800 3056 197245 3336
rect 800 2384 197695 3056
rect 880 2143 197695 2384
<< metal4 >>
rect 4208 2128 4528 198064
rect 19568 2128 19888 198064
rect 34928 2128 35248 198064
rect 50288 2128 50608 198064
rect 65648 2128 65968 198064
rect 81008 2128 81328 198064
rect 96368 2128 96688 198064
rect 111728 2128 112048 198064
rect 127088 2128 127408 198064
rect 142448 2128 142768 198064
rect 157808 2128 158128 198064
rect 173168 2128 173488 198064
rect 188528 2128 188848 198064
<< obsm4 >>
rect 10915 198144 195533 198389
rect 10915 2891 19488 198144
rect 19968 2891 34848 198144
rect 35328 2891 50208 198144
rect 50688 2891 65568 198144
rect 66048 2891 80928 198144
rect 81408 2891 96288 198144
rect 96768 2891 111648 198144
rect 112128 2891 127008 198144
rect 127488 2891 142368 198144
rect 142848 2891 157728 198144
rect 158208 2891 173088 198144
rect 173568 2891 188448 198144
rect 188928 2891 195533 198144
<< labels >>
rlabel metal3 s 197325 3136 198125 3256 6 clk_i
port 1 nsew signal input
rlabel metal2 s 146298 199469 146354 200269 6 i_dout0[0]
port 2 nsew signal input
rlabel metal2 s 163778 0 163834 800 6 i_dout0[10]
port 3 nsew signal input
rlabel metal2 s 166446 0 166502 800 6 i_dout0[11]
port 4 nsew signal input
rlabel metal2 s 169022 0 169078 800 6 i_dout0[12]
port 5 nsew signal input
rlabel metal3 s 197325 99968 198125 100088 6 i_dout0[13]
port 6 nsew signal input
rlabel metal3 s 0 115880 800 116000 6 i_dout0[14]
port 7 nsew signal input
rlabel metal3 s 0 120504 800 120624 6 i_dout0[15]
port 8 nsew signal input
rlabel metal2 s 176934 199469 176990 200269 6 i_dout0[16]
port 9 nsew signal input
rlabel metal2 s 175462 0 175518 800 6 i_dout0[17]
port 10 nsew signal input
rlabel metal2 s 179510 199469 179566 200269 6 i_dout0[18]
port 11 nsew signal input
rlabel metal2 s 178038 0 178094 800 6 i_dout0[19]
port 12 nsew signal input
rlabel metal3 s 197325 28976 198125 29096 6 i_dout0[1]
port 13 nsew signal input
rlabel metal2 s 180798 199469 180854 200269 6 i_dout0[20]
port 14 nsew signal input
rlabel metal2 s 179326 0 179382 800 6 i_dout0[21]
port 15 nsew signal input
rlabel metal3 s 0 170552 800 170672 6 i_dout0[22]
port 16 nsew signal input
rlabel metal3 s 0 175176 800 175296 6 i_dout0[23]
port 17 nsew signal input
rlabel metal3 s 0 179664 800 179784 6 i_dout0[24]
port 18 nsew signal input
rlabel metal3 s 0 184288 800 184408 6 i_dout0[25]
port 19 nsew signal input
rlabel metal2 s 193586 199469 193642 200269 6 i_dout0[26]
port 20 nsew signal input
rlabel metal2 s 184570 0 184626 800 6 i_dout0[27]
port 21 nsew signal input
rlabel metal3 s 197325 184016 198125 184136 6 i_dout0[28]
port 22 nsew signal input
rlabel metal2 s 196162 199469 196218 200269 6 i_dout0[29]
port 23 nsew signal input
rlabel metal3 s 0 43120 800 43240 6 i_dout0[2]
port 24 nsew signal input
rlabel metal2 s 192298 0 192354 800 6 i_dout0[30]
port 25 nsew signal input
rlabel metal3 s 197325 196936 198125 197056 6 i_dout0[31]
port 26 nsew signal input
rlabel metal3 s 0 47608 800 47728 6 i_dout0[3]
port 27 nsew signal input
rlabel metal3 s 0 61344 800 61464 6 i_dout0[4]
port 28 nsew signal input
rlabel metal2 s 153474 0 153530 800 6 i_dout0[5]
port 29 nsew signal input
rlabel metal3 s 197325 67736 198125 67856 6 i_dout0[6]
port 30 nsew signal input
rlabel metal2 s 164146 199469 164202 200269 6 i_dout0[7]
port 31 nsew signal input
rlabel metal3 s 0 88680 800 88800 6 i_dout0[8]
port 32 nsew signal input
rlabel metal3 s 0 102280 800 102400 6 i_dout0[9]
port 33 nsew signal input
rlabel metal3 s 0 11160 800 11280 6 i_dout0_1[0]
port 34 nsew signal input
rlabel metal2 s 170586 199469 170642 200269 6 i_dout0_1[10]
port 35 nsew signal input
rlabel metal2 s 165066 0 165122 800 6 i_dout0_1[11]
port 36 nsew signal input
rlabel metal2 s 167734 0 167790 800 6 i_dout0_1[12]
port 37 nsew signal input
rlabel metal3 s 0 106768 800 106888 6 i_dout0_1[13]
port 38 nsew signal input
rlabel metal3 s 197325 106496 198125 106616 6 i_dout0_1[14]
port 39 nsew signal input
rlabel metal2 s 175646 199469 175702 200269 6 i_dout0_1[15]
port 40 nsew signal input
rlabel metal3 s 0 124992 800 125112 6 i_dout0_1[16]
port 41 nsew signal input
rlabel metal3 s 0 129616 800 129736 6 i_dout0_1[17]
port 42 nsew signal input
rlabel metal3 s 197325 132336 198125 132456 6 i_dout0_1[18]
port 43 nsew signal input
rlabel metal3 s 0 147840 800 147960 6 i_dout0_1[19]
port 44 nsew signal input
rlabel metal3 s 0 29384 800 29504 6 i_dout0_1[1]
port 45 nsew signal input
rlabel metal3 s 197325 145256 198125 145376 6 i_dout0_1[20]
port 46 nsew signal input
rlabel metal3 s 0 161440 800 161560 6 i_dout0_1[21]
port 47 nsew signal input
rlabel metal2 s 183374 199469 183430 200269 6 i_dout0_1[22]
port 48 nsew signal input
rlabel metal2 s 184662 199469 184718 200269 6 i_dout0_1[23]
port 49 nsew signal input
rlabel metal2 s 180614 0 180670 800 6 i_dout0_1[24]
port 50 nsew signal input
rlabel metal2 s 189722 199469 189778 200269 6 i_dout0_1[25]
port 51 nsew signal input
rlabel metal3 s 0 188776 800 188896 6 i_dout0_1[26]
port 52 nsew signal input
rlabel metal2 s 183282 0 183338 800 6 i_dout0_1[27]
port 53 nsew signal input
rlabel metal2 s 187146 0 187202 800 6 i_dout0_1[28]
port 54 nsew signal input
rlabel metal2 s 194874 199469 194930 200269 6 i_dout0_1[29]
port 55 nsew signal input
rlabel metal3 s 197325 41896 198125 42016 6 i_dout0_1[2]
port 56 nsew signal input
rlabel metal2 s 191010 0 191066 800 6 i_dout0_1[30]
port 57 nsew signal input
rlabel metal2 s 196162 0 196218 800 6 i_dout0_1[31]
port 58 nsew signal input
rlabel metal2 s 149610 0 149666 800 6 i_dout0_1[3]
port 59 nsew signal input
rlabel metal3 s 197325 61208 198125 61328 6 i_dout0_1[4]
port 60 nsew signal input
rlabel metal2 s 159086 199469 159142 200269 6 i_dout0_1[5]
port 61 nsew signal input
rlabel metal3 s 0 79568 800 79688 6 i_dout0_1[6]
port 62 nsew signal input
rlabel metal2 s 157338 0 157394 800 6 i_dout0_1[7]
port 63 nsew signal input
rlabel metal2 s 161202 0 161258 800 6 i_dout0_1[8]
port 64 nsew signal input
rlabel metal2 s 168010 199469 168066 200269 6 i_dout0_1[9]
port 65 nsew signal input
rlabel metal2 s 570 199469 626 200269 6 io_in[0]
port 66 nsew signal input
rlabel metal2 s 38842 199469 38898 200269 6 io_in[10]
port 67 nsew signal input
rlabel metal2 s 42706 199469 42762 200269 6 io_in[11]
port 68 nsew signal input
rlabel metal2 s 46570 199469 46626 200269 6 io_in[12]
port 69 nsew signal input
rlabel metal2 s 50342 199469 50398 200269 6 io_in[13]
port 70 nsew signal input
rlabel metal2 s 54206 199469 54262 200269 6 io_in[14]
port 71 nsew signal input
rlabel metal2 s 58070 199469 58126 200269 6 io_in[15]
port 72 nsew signal input
rlabel metal2 s 61934 199469 61990 200269 6 io_in[16]
port 73 nsew signal input
rlabel metal2 s 65706 199469 65762 200269 6 io_in[17]
port 74 nsew signal input
rlabel metal2 s 69570 199469 69626 200269 6 io_in[18]
port 75 nsew signal input
rlabel metal2 s 73434 199469 73490 200269 6 io_in[19]
port 76 nsew signal input
rlabel metal2 s 4342 199469 4398 200269 6 io_in[1]
port 77 nsew signal input
rlabel metal2 s 77206 199469 77262 200269 6 io_in[20]
port 78 nsew signal input
rlabel metal2 s 81070 199469 81126 200269 6 io_in[21]
port 79 nsew signal input
rlabel metal2 s 84934 199469 84990 200269 6 io_in[22]
port 80 nsew signal input
rlabel metal2 s 88706 199469 88762 200269 6 io_in[23]
port 81 nsew signal input
rlabel metal2 s 92570 199469 92626 200269 6 io_in[24]
port 82 nsew signal input
rlabel metal2 s 96434 199469 96490 200269 6 io_in[25]
port 83 nsew signal input
rlabel metal2 s 100206 199469 100262 200269 6 io_in[26]
port 84 nsew signal input
rlabel metal2 s 104070 199469 104126 200269 6 io_in[27]
port 85 nsew signal input
rlabel metal2 s 107934 199469 107990 200269 6 io_in[28]
port 86 nsew signal input
rlabel metal2 s 111798 199469 111854 200269 6 io_in[29]
port 87 nsew signal input
rlabel metal2 s 8206 199469 8262 200269 6 io_in[2]
port 88 nsew signal input
rlabel metal2 s 115570 199469 115626 200269 6 io_in[30]
port 89 nsew signal input
rlabel metal2 s 119434 199469 119490 200269 6 io_in[31]
port 90 nsew signal input
rlabel metal2 s 123298 199469 123354 200269 6 io_in[32]
port 91 nsew signal input
rlabel metal2 s 127070 199469 127126 200269 6 io_in[33]
port 92 nsew signal input
rlabel metal2 s 130934 199469 130990 200269 6 io_in[34]
port 93 nsew signal input
rlabel metal2 s 134798 199469 134854 200269 6 io_in[35]
port 94 nsew signal input
rlabel metal2 s 138570 199469 138626 200269 6 io_in[36]
port 95 nsew signal input
rlabel metal2 s 142434 199469 142490 200269 6 io_in[37]
port 96 nsew signal input
rlabel metal2 s 12070 199469 12126 200269 6 io_in[3]
port 97 nsew signal input
rlabel metal2 s 15842 199469 15898 200269 6 io_in[4]
port 98 nsew signal input
rlabel metal2 s 19706 199469 19762 200269 6 io_in[5]
port 99 nsew signal input
rlabel metal2 s 23570 199469 23626 200269 6 io_in[6]
port 100 nsew signal input
rlabel metal2 s 27342 199469 27398 200269 6 io_in[7]
port 101 nsew signal input
rlabel metal2 s 31206 199469 31262 200269 6 io_in[8]
port 102 nsew signal input
rlabel metal2 s 35070 199469 35126 200269 6 io_in[9]
port 103 nsew signal input
rlabel metal2 s 1766 199469 1822 200269 6 io_oeb[0]
port 104 nsew signal output
rlabel metal2 s 40130 199469 40186 200269 6 io_oeb[10]
port 105 nsew signal output
rlabel metal2 s 43994 199469 44050 200269 6 io_oeb[11]
port 106 nsew signal output
rlabel metal2 s 47858 199469 47914 200269 6 io_oeb[12]
port 107 nsew signal output
rlabel metal2 s 51630 199469 51686 200269 6 io_oeb[13]
port 108 nsew signal output
rlabel metal2 s 55494 199469 55550 200269 6 io_oeb[14]
port 109 nsew signal output
rlabel metal2 s 59358 199469 59414 200269 6 io_oeb[15]
port 110 nsew signal output
rlabel metal2 s 63130 199469 63186 200269 6 io_oeb[16]
port 111 nsew signal output
rlabel metal2 s 66994 199469 67050 200269 6 io_oeb[17]
port 112 nsew signal output
rlabel metal2 s 70858 199469 70914 200269 6 io_oeb[18]
port 113 nsew signal output
rlabel metal2 s 74722 199469 74778 200269 6 io_oeb[19]
port 114 nsew signal output
rlabel metal2 s 5630 199469 5686 200269 6 io_oeb[1]
port 115 nsew signal output
rlabel metal2 s 78494 199469 78550 200269 6 io_oeb[20]
port 116 nsew signal output
rlabel metal2 s 82358 199469 82414 200269 6 io_oeb[21]
port 117 nsew signal output
rlabel metal2 s 86222 199469 86278 200269 6 io_oeb[22]
port 118 nsew signal output
rlabel metal2 s 89994 199469 90050 200269 6 io_oeb[23]
port 119 nsew signal output
rlabel metal2 s 93858 199469 93914 200269 6 io_oeb[24]
port 120 nsew signal output
rlabel metal2 s 97722 199469 97778 200269 6 io_oeb[25]
port 121 nsew signal output
rlabel metal2 s 101494 199469 101550 200269 6 io_oeb[26]
port 122 nsew signal output
rlabel metal2 s 105358 199469 105414 200269 6 io_oeb[27]
port 123 nsew signal output
rlabel metal2 s 109222 199469 109278 200269 6 io_oeb[28]
port 124 nsew signal output
rlabel metal2 s 112994 199469 113050 200269 6 io_oeb[29]
port 125 nsew signal output
rlabel metal2 s 9494 199469 9550 200269 6 io_oeb[2]
port 126 nsew signal output
rlabel metal2 s 116858 199469 116914 200269 6 io_oeb[30]
port 127 nsew signal output
rlabel metal2 s 120722 199469 120778 200269 6 io_oeb[31]
port 128 nsew signal output
rlabel metal2 s 124494 199469 124550 200269 6 io_oeb[32]
port 129 nsew signal output
rlabel metal2 s 128358 199469 128414 200269 6 io_oeb[33]
port 130 nsew signal output
rlabel metal2 s 132222 199469 132278 200269 6 io_oeb[34]
port 131 nsew signal output
rlabel metal2 s 136086 199469 136142 200269 6 io_oeb[35]
port 132 nsew signal output
rlabel metal2 s 139858 199469 139914 200269 6 io_oeb[36]
port 133 nsew signal output
rlabel metal2 s 143722 199469 143778 200269 6 io_oeb[37]
port 134 nsew signal output
rlabel metal2 s 13266 199469 13322 200269 6 io_oeb[3]
port 135 nsew signal output
rlabel metal2 s 17130 199469 17186 200269 6 io_oeb[4]
port 136 nsew signal output
rlabel metal2 s 20994 199469 21050 200269 6 io_oeb[5]
port 137 nsew signal output
rlabel metal2 s 24858 199469 24914 200269 6 io_oeb[6]
port 138 nsew signal output
rlabel metal2 s 28630 199469 28686 200269 6 io_oeb[7]
port 139 nsew signal output
rlabel metal2 s 32494 199469 32550 200269 6 io_oeb[8]
port 140 nsew signal output
rlabel metal2 s 36358 199469 36414 200269 6 io_oeb[9]
port 141 nsew signal output
rlabel metal2 s 3054 199469 3110 200269 6 io_out[0]
port 142 nsew signal output
rlabel metal2 s 41418 199469 41474 200269 6 io_out[10]
port 143 nsew signal output
rlabel metal2 s 45282 199469 45338 200269 6 io_out[11]
port 144 nsew signal output
rlabel metal2 s 49146 199469 49202 200269 6 io_out[12]
port 145 nsew signal output
rlabel metal2 s 52918 199469 52974 200269 6 io_out[13]
port 146 nsew signal output
rlabel metal2 s 56782 199469 56838 200269 6 io_out[14]
port 147 nsew signal output
rlabel metal2 s 60646 199469 60702 200269 6 io_out[15]
port 148 nsew signal output
rlabel metal2 s 64418 199469 64474 200269 6 io_out[16]
port 149 nsew signal output
rlabel metal2 s 68282 199469 68338 200269 6 io_out[17]
port 150 nsew signal output
rlabel metal2 s 72146 199469 72202 200269 6 io_out[18]
port 151 nsew signal output
rlabel metal2 s 75918 199469 75974 200269 6 io_out[19]
port 152 nsew signal output
rlabel metal2 s 6918 199469 6974 200269 6 io_out[1]
port 153 nsew signal output
rlabel metal2 s 79782 199469 79838 200269 6 io_out[20]
port 154 nsew signal output
rlabel metal2 s 83646 199469 83702 200269 6 io_out[21]
port 155 nsew signal output
rlabel metal2 s 87418 199469 87474 200269 6 io_out[22]
port 156 nsew signal output
rlabel metal2 s 91282 199469 91338 200269 6 io_out[23]
port 157 nsew signal output
rlabel metal2 s 95146 199469 95202 200269 6 io_out[24]
port 158 nsew signal output
rlabel metal2 s 99010 199469 99066 200269 6 io_out[25]
port 159 nsew signal output
rlabel metal2 s 102782 199469 102838 200269 6 io_out[26]
port 160 nsew signal output
rlabel metal2 s 106646 199469 106702 200269 6 io_out[27]
port 161 nsew signal output
rlabel metal2 s 110510 199469 110566 200269 6 io_out[28]
port 162 nsew signal output
rlabel metal2 s 114282 199469 114338 200269 6 io_out[29]
port 163 nsew signal output
rlabel metal2 s 10782 199469 10838 200269 6 io_out[2]
port 164 nsew signal output
rlabel metal2 s 118146 199469 118202 200269 6 io_out[30]
port 165 nsew signal output
rlabel metal2 s 122010 199469 122066 200269 6 io_out[31]
port 166 nsew signal output
rlabel metal2 s 125782 199469 125838 200269 6 io_out[32]
port 167 nsew signal output
rlabel metal2 s 129646 199469 129702 200269 6 io_out[33]
port 168 nsew signal output
rlabel metal2 s 133510 199469 133566 200269 6 io_out[34]
port 169 nsew signal output
rlabel metal2 s 137282 199469 137338 200269 6 io_out[35]
port 170 nsew signal output
rlabel metal2 s 141146 199469 141202 200269 6 io_out[36]
port 171 nsew signal output
rlabel metal2 s 145010 199469 145066 200269 6 io_out[37]
port 172 nsew signal output
rlabel metal2 s 14554 199469 14610 200269 6 io_out[3]
port 173 nsew signal output
rlabel metal2 s 18418 199469 18474 200269 6 io_out[4]
port 174 nsew signal output
rlabel metal2 s 22282 199469 22338 200269 6 io_out[5]
port 175 nsew signal output
rlabel metal2 s 26054 199469 26110 200269 6 io_out[6]
port 176 nsew signal output
rlabel metal2 s 29918 199469 29974 200269 6 io_out[7]
port 177 nsew signal output
rlabel metal2 s 33782 199469 33838 200269 6 io_out[8]
port 178 nsew signal output
rlabel metal2 s 37646 199469 37702 200269 6 io_out[9]
port 179 nsew signal output
rlabel metal2 s 137926 0 137982 800 6 irq[0]
port 180 nsew signal output
rlabel metal2 s 139214 0 139270 800 6 irq[1]
port 181 nsew signal output
rlabel metal2 s 140502 0 140558 800 6 irq[2]
port 182 nsew signal output
rlabel metal3 s 0 2184 800 2304 6 o_csb0
port 183 nsew signal output
rlabel metal3 s 197325 9528 198125 9648 6 o_csb0_1
port 184 nsew signal output
rlabel metal2 s 147586 199469 147642 200269 6 o_din0[0]
port 185 nsew signal output
rlabel metal2 s 173162 199469 173218 200269 6 o_din0[10]
port 186 nsew signal output
rlabel metal3 s 197325 93576 198125 93696 6 o_din0[11]
port 187 nsew signal output
rlabel metal2 s 171598 0 171654 800 6 o_din0[12]
port 188 nsew signal output
rlabel metal3 s 0 111392 800 111512 6 o_din0[13]
port 189 nsew signal output
rlabel metal2 s 174174 0 174230 800 6 o_din0[14]
port 190 nsew signal output
rlabel metal3 s 197325 119416 198125 119536 6 o_din0[15]
port 191 nsew signal output
rlabel metal3 s 197325 125808 198125 125928 6 o_din0[16]
port 192 nsew signal output
rlabel metal3 s 0 134104 800 134224 6 o_din0[17]
port 193 nsew signal output
rlabel metal3 s 0 143216 800 143336 6 o_din0[18]
port 194 nsew signal output
rlabel metal3 s 0 152328 800 152448 6 o_din0[19]
port 195 nsew signal output
rlabel metal2 s 150070 199469 150126 200269 6 o_din0[1]
port 196 nsew signal output
rlabel metal3 s 0 156952 800 157072 6 o_din0[20]
port 197 nsew signal output
rlabel metal3 s 0 166064 800 166184 6 o_din0[21]
port 198 nsew signal output
rlabel metal3 s 197325 164568 198125 164688 6 o_din0[22]
port 199 nsew signal output
rlabel metal2 s 185950 199469 186006 200269 6 o_din0[23]
port 200 nsew signal output
rlabel metal2 s 188434 199469 188490 200269 6 o_din0[24]
port 201 nsew signal output
rlabel metal2 s 192298 199469 192354 200269 6 o_din0[25]
port 202 nsew signal output
rlabel metal3 s 0 193400 800 193520 6 o_din0[26]
port 203 nsew signal output
rlabel metal2 s 185858 0 185914 800 6 o_din0[27]
port 204 nsew signal output
rlabel metal3 s 0 197888 800 198008 6 o_din0[28]
port 205 nsew signal output
rlabel metal3 s 197325 190408 198125 190528 6 o_din0[29]
port 206 nsew signal output
rlabel metal2 s 145654 0 145710 800 6 o_din0[2]
port 207 nsew signal output
rlabel metal2 s 194874 0 194930 800 6 o_din0[30]
port 208 nsew signal output
rlabel metal2 s 197450 0 197506 800 6 o_din0[31]
port 209 nsew signal output
rlabel metal3 s 197325 54816 198125 54936 6 o_din0[3]
port 210 nsew signal output
rlabel metal3 s 0 65832 800 65952 6 o_din0[4]
port 211 nsew signal output
rlabel metal3 s 0 70456 800 70576 6 o_din0[5]
port 212 nsew signal output
rlabel metal2 s 162858 199469 162914 200269 6 o_din0[6]
port 213 nsew signal output
rlabel metal3 s 0 84056 800 84176 6 o_din0[7]
port 214 nsew signal output
rlabel metal3 s 0 93168 800 93288 6 o_din0[8]
port 215 nsew signal output
rlabel metal2 s 162490 0 162546 800 6 o_din0[9]
port 216 nsew signal output
rlabel metal2 s 148874 199469 148930 200269 6 o_din0_1[0]
port 217 nsew signal output
rlabel metal2 s 171874 199469 171930 200269 6 o_din0_1[10]
port 218 nsew signal output
rlabel metal3 s 197325 87048 198125 87168 6 o_din0_1[11]
port 219 nsew signal output
rlabel metal2 s 170310 0 170366 800 6 o_din0_1[12]
port 220 nsew signal output
rlabel metal2 s 174358 199469 174414 200269 6 o_din0_1[13]
port 221 nsew signal output
rlabel metal2 s 172886 0 172942 800 6 o_din0_1[14]
port 222 nsew signal output
rlabel metal3 s 197325 112888 198125 113008 6 o_din0_1[15]
port 223 nsew signal output
rlabel metal2 s 178222 199469 178278 200269 6 o_din0_1[16]
port 224 nsew signal output
rlabel metal2 s 176750 0 176806 800 6 o_din0_1[17]
port 225 nsew signal output
rlabel metal3 s 0 138728 800 138848 6 o_din0_1[18]
port 226 nsew signal output
rlabel metal3 s 197325 138728 198125 138848 6 o_din0_1[19]
port 227 nsew signal output
rlabel metal3 s 197325 35368 198125 35488 6 o_din0_1[1]
port 228 nsew signal output
rlabel metal2 s 182086 199469 182142 200269 6 o_din0_1[20]
port 229 nsew signal output
rlabel metal3 s 197325 151648 198125 151768 6 o_din0_1[21]
port 230 nsew signal output
rlabel metal3 s 197325 158176 198125 158296 6 o_din0_1[22]
port 231 nsew signal output
rlabel metal3 s 197325 171096 198125 171216 6 o_din0_1[23]
port 232 nsew signal output
rlabel metal2 s 187146 199469 187202 200269 6 o_din0_1[24]
port 233 nsew signal output
rlabel metal2 s 191010 199469 191066 200269 6 o_din0_1[25]
port 234 nsew signal output
rlabel metal2 s 181902 0 181958 800 6 o_din0_1[26]
port 235 nsew signal output
rlabel metal3 s 197325 177488 198125 177608 6 o_din0_1[27]
port 236 nsew signal output
rlabel metal2 s 188434 0 188490 800 6 o_din0_1[28]
port 237 nsew signal output
rlabel metal2 s 189722 0 189778 800 6 o_din0_1[29]
port 238 nsew signal output
rlabel metal3 s 197325 48288 198125 48408 6 o_din0_1[2]
port 239 nsew signal output
rlabel metal2 s 193586 0 193642 800 6 o_din0_1[30]
port 240 nsew signal output
rlabel metal2 s 197450 199469 197506 200269 6 o_din0_1[31]
port 241 nsew signal output
rlabel metal2 s 153934 199469 153990 200269 6 o_din0_1[3]
port 242 nsew signal output
rlabel metal2 s 155222 199469 155278 200269 6 o_din0_1[4]
port 243 nsew signal output
rlabel metal2 s 160374 199469 160430 200269 6 o_din0_1[5]
port 244 nsew signal output
rlabel metal2 s 161570 199469 161626 200269 6 o_din0_1[6]
port 245 nsew signal output
rlabel metal2 s 158626 0 158682 800 6 o_din0_1[7]
port 246 nsew signal output
rlabel metal3 s 197325 80656 198125 80776 6 o_din0_1[8]
port 247 nsew signal output
rlabel metal2 s 169298 199469 169354 200269 6 o_din0_1[9]
port 248 nsew signal output
rlabel metal3 s 0 15784 800 15904 6 o_waddr0[0]
port 249 nsew signal output
rlabel metal2 s 144366 0 144422 800 6 o_waddr0[1]
port 250 nsew signal output
rlabel metal2 s 152646 199469 152702 200269 6 o_waddr0[2]
port 251 nsew signal output
rlabel metal2 s 150898 0 150954 800 6 o_waddr0[3]
port 252 nsew signal output
rlabel metal2 s 157798 199469 157854 200269 6 o_waddr0[4]
port 253 nsew signal output
rlabel metal2 s 154762 0 154818 800 6 o_waddr0[5]
port 254 nsew signal output
rlabel metal3 s 197325 74128 198125 74248 6 o_waddr0[6]
port 255 nsew signal output
rlabel metal2 s 159914 0 159970 800 6 o_waddr0[7]
port 256 nsew signal output
rlabel metal3 s 0 97792 800 97912 6 o_waddr0[8]
port 257 nsew signal output
rlabel metal3 s 0 20272 800 20392 6 o_waddr0_1[0]
port 258 nsew signal output
rlabel metal2 s 143078 0 143134 800 6 o_waddr0_1[1]
port 259 nsew signal output
rlabel metal2 s 151358 199469 151414 200269 6 o_waddr0_1[2]
port 260 nsew signal output
rlabel metal3 s 0 52232 800 52352 6 o_waddr0_1[3]
port 261 nsew signal output
rlabel metal2 s 156510 199469 156566 200269 6 o_waddr0_1[4]
port 262 nsew signal output
rlabel metal3 s 0 74944 800 75064 6 o_waddr0_1[5]
port 263 nsew signal output
rlabel metal2 s 156050 0 156106 800 6 o_waddr0_1[6]
port 264 nsew signal output
rlabel metal2 s 165434 199469 165490 200269 6 o_waddr0_1[7]
port 265 nsew signal output
rlabel metal2 s 166722 199469 166778 200269 6 o_waddr0_1[8]
port 266 nsew signal output
rlabel metal3 s 0 6672 800 6792 6 o_web0
port 267 nsew signal output
rlabel metal3 s 197325 16056 198125 16176 6 o_web0_1
port 268 nsew signal output
rlabel metal2 s 141790 0 141846 800 6 o_wmask0[0]
port 269 nsew signal output
rlabel metal3 s 0 38496 800 38616 6 o_wmask0[1]
port 270 nsew signal output
rlabel metal2 s 148230 0 148286 800 6 o_wmask0[2]
port 271 nsew signal output
rlabel metal3 s 0 56720 800 56840 6 o_wmask0[3]
port 272 nsew signal output
rlabel metal3 s 0 24896 800 25016 6 o_wmask0_1[0]
port 273 nsew signal output
rlabel metal3 s 0 34008 800 34128 6 o_wmask0_1[1]
port 274 nsew signal output
rlabel metal2 s 146942 0 146998 800 6 o_wmask0_1[2]
port 275 nsew signal output
rlabel metal2 s 152186 0 152242 800 6 o_wmask0_1[3]
port 276 nsew signal output
rlabel metal3 s 197325 22448 198125 22568 6 rst_i
port 277 nsew signal input
rlabel metal4 s 4208 2128 4528 198064 6 vccd1
port 278 nsew power input
rlabel metal4 s 34928 2128 35248 198064 6 vccd1
port 278 nsew power input
rlabel metal4 s 65648 2128 65968 198064 6 vccd1
port 278 nsew power input
rlabel metal4 s 96368 2128 96688 198064 6 vccd1
port 278 nsew power input
rlabel metal4 s 127088 2128 127408 198064 6 vccd1
port 278 nsew power input
rlabel metal4 s 157808 2128 158128 198064 6 vccd1
port 278 nsew power input
rlabel metal4 s 188528 2128 188848 198064 6 vccd1
port 278 nsew power input
rlabel metal4 s 19568 2128 19888 198064 6 vssd1
port 279 nsew ground input
rlabel metal4 s 50288 2128 50608 198064 6 vssd1
port 279 nsew ground input
rlabel metal4 s 81008 2128 81328 198064 6 vssd1
port 279 nsew ground input
rlabel metal4 s 111728 2128 112048 198064 6 vssd1
port 279 nsew ground input
rlabel metal4 s 142448 2128 142768 198064 6 vssd1
port 279 nsew ground input
rlabel metal4 s 173168 2128 173488 198064 6 vssd1
port 279 nsew ground input
rlabel metal2 s 662 0 718 800 6 wb_clk_i
port 280 nsew signal input
rlabel metal2 s 1950 0 2006 800 6 wb_rst_i
port 281 nsew signal input
rlabel metal2 s 3238 0 3294 800 6 wbs_ack_o
port 282 nsew signal output
rlabel metal2 s 8390 0 8446 800 6 wbs_adr_i[0]
port 283 nsew signal input
rlabel metal2 s 52458 0 52514 800 6 wbs_adr_i[10]
port 284 nsew signal input
rlabel metal2 s 56322 0 56378 800 6 wbs_adr_i[11]
port 285 nsew signal input
rlabel metal2 s 60186 0 60242 800 6 wbs_adr_i[12]
port 286 nsew signal input
rlabel metal2 s 64050 0 64106 800 6 wbs_adr_i[13]
port 287 nsew signal input
rlabel metal2 s 68006 0 68062 800 6 wbs_adr_i[14]
port 288 nsew signal input
rlabel metal2 s 71870 0 71926 800 6 wbs_adr_i[15]
port 289 nsew signal input
rlabel metal2 s 75734 0 75790 800 6 wbs_adr_i[16]
port 290 nsew signal input
rlabel metal2 s 79598 0 79654 800 6 wbs_adr_i[17]
port 291 nsew signal input
rlabel metal2 s 83554 0 83610 800 6 wbs_adr_i[18]
port 292 nsew signal input
rlabel metal2 s 87418 0 87474 800 6 wbs_adr_i[19]
port 293 nsew signal input
rlabel metal2 s 13542 0 13598 800 6 wbs_adr_i[1]
port 294 nsew signal input
rlabel metal2 s 91282 0 91338 800 6 wbs_adr_i[20]
port 295 nsew signal input
rlabel metal2 s 95146 0 95202 800 6 wbs_adr_i[21]
port 296 nsew signal input
rlabel metal2 s 99010 0 99066 800 6 wbs_adr_i[22]
port 297 nsew signal input
rlabel metal2 s 102966 0 103022 800 6 wbs_adr_i[23]
port 298 nsew signal input
rlabel metal2 s 106830 0 106886 800 6 wbs_adr_i[24]
port 299 nsew signal input
rlabel metal2 s 110694 0 110750 800 6 wbs_adr_i[25]
port 300 nsew signal input
rlabel metal2 s 114558 0 114614 800 6 wbs_adr_i[26]
port 301 nsew signal input
rlabel metal2 s 118514 0 118570 800 6 wbs_adr_i[27]
port 302 nsew signal input
rlabel metal2 s 122378 0 122434 800 6 wbs_adr_i[28]
port 303 nsew signal input
rlabel metal2 s 126242 0 126298 800 6 wbs_adr_i[29]
port 304 nsew signal input
rlabel metal2 s 18786 0 18842 800 6 wbs_adr_i[2]
port 305 nsew signal input
rlabel metal2 s 130106 0 130162 800 6 wbs_adr_i[30]
port 306 nsew signal input
rlabel metal2 s 134062 0 134118 800 6 wbs_adr_i[31]
port 307 nsew signal input
rlabel metal2 s 23938 0 23994 800 6 wbs_adr_i[3]
port 308 nsew signal input
rlabel metal2 s 29090 0 29146 800 6 wbs_adr_i[4]
port 309 nsew signal input
rlabel metal2 s 32954 0 33010 800 6 wbs_adr_i[5]
port 310 nsew signal input
rlabel metal2 s 36910 0 36966 800 6 wbs_adr_i[6]
port 311 nsew signal input
rlabel metal2 s 40774 0 40830 800 6 wbs_adr_i[7]
port 312 nsew signal input
rlabel metal2 s 44638 0 44694 800 6 wbs_adr_i[8]
port 313 nsew signal input
rlabel metal2 s 48502 0 48558 800 6 wbs_adr_i[9]
port 314 nsew signal input
rlabel metal2 s 4526 0 4582 800 6 wbs_cyc_i
port 315 nsew signal input
rlabel metal2 s 9678 0 9734 800 6 wbs_dat_i[0]
port 316 nsew signal input
rlabel metal2 s 53746 0 53802 800 6 wbs_dat_i[10]
port 317 nsew signal input
rlabel metal2 s 57610 0 57666 800 6 wbs_dat_i[11]
port 318 nsew signal input
rlabel metal2 s 61474 0 61530 800 6 wbs_dat_i[12]
port 319 nsew signal input
rlabel metal2 s 65338 0 65394 800 6 wbs_dat_i[13]
port 320 nsew signal input
rlabel metal2 s 69294 0 69350 800 6 wbs_dat_i[14]
port 321 nsew signal input
rlabel metal2 s 73158 0 73214 800 6 wbs_dat_i[15]
port 322 nsew signal input
rlabel metal2 s 77022 0 77078 800 6 wbs_dat_i[16]
port 323 nsew signal input
rlabel metal2 s 80886 0 80942 800 6 wbs_dat_i[17]
port 324 nsew signal input
rlabel metal2 s 84842 0 84898 800 6 wbs_dat_i[18]
port 325 nsew signal input
rlabel metal2 s 88706 0 88762 800 6 wbs_dat_i[19]
port 326 nsew signal input
rlabel metal2 s 14830 0 14886 800 6 wbs_dat_i[1]
port 327 nsew signal input
rlabel metal2 s 92570 0 92626 800 6 wbs_dat_i[20]
port 328 nsew signal input
rlabel metal2 s 96434 0 96490 800 6 wbs_dat_i[21]
port 329 nsew signal input
rlabel metal2 s 100390 0 100446 800 6 wbs_dat_i[22]
port 330 nsew signal input
rlabel metal2 s 104254 0 104310 800 6 wbs_dat_i[23]
port 331 nsew signal input
rlabel metal2 s 108118 0 108174 800 6 wbs_dat_i[24]
port 332 nsew signal input
rlabel metal2 s 111982 0 112038 800 6 wbs_dat_i[25]
port 333 nsew signal input
rlabel metal2 s 115846 0 115902 800 6 wbs_dat_i[26]
port 334 nsew signal input
rlabel metal2 s 119802 0 119858 800 6 wbs_dat_i[27]
port 335 nsew signal input
rlabel metal2 s 123666 0 123722 800 6 wbs_dat_i[28]
port 336 nsew signal input
rlabel metal2 s 127530 0 127586 800 6 wbs_dat_i[29]
port 337 nsew signal input
rlabel metal2 s 20074 0 20130 800 6 wbs_dat_i[2]
port 338 nsew signal input
rlabel metal2 s 131394 0 131450 800 6 wbs_dat_i[30]
port 339 nsew signal input
rlabel metal2 s 135350 0 135406 800 6 wbs_dat_i[31]
port 340 nsew signal input
rlabel metal2 s 25226 0 25282 800 6 wbs_dat_i[3]
port 341 nsew signal input
rlabel metal2 s 30378 0 30434 800 6 wbs_dat_i[4]
port 342 nsew signal input
rlabel metal2 s 34334 0 34390 800 6 wbs_dat_i[5]
port 343 nsew signal input
rlabel metal2 s 38198 0 38254 800 6 wbs_dat_i[6]
port 344 nsew signal input
rlabel metal2 s 42062 0 42118 800 6 wbs_dat_i[7]
port 345 nsew signal input
rlabel metal2 s 45926 0 45982 800 6 wbs_dat_i[8]
port 346 nsew signal input
rlabel metal2 s 49790 0 49846 800 6 wbs_dat_i[9]
port 347 nsew signal input
rlabel metal2 s 10966 0 11022 800 6 wbs_dat_o[0]
port 348 nsew signal output
rlabel metal2 s 55034 0 55090 800 6 wbs_dat_o[10]
port 349 nsew signal output
rlabel metal2 s 58898 0 58954 800 6 wbs_dat_o[11]
port 350 nsew signal output
rlabel metal2 s 62762 0 62818 800 6 wbs_dat_o[12]
port 351 nsew signal output
rlabel metal2 s 66718 0 66774 800 6 wbs_dat_o[13]
port 352 nsew signal output
rlabel metal2 s 70582 0 70638 800 6 wbs_dat_o[14]
port 353 nsew signal output
rlabel metal2 s 74446 0 74502 800 6 wbs_dat_o[15]
port 354 nsew signal output
rlabel metal2 s 78310 0 78366 800 6 wbs_dat_o[16]
port 355 nsew signal output
rlabel metal2 s 82174 0 82230 800 6 wbs_dat_o[17]
port 356 nsew signal output
rlabel metal2 s 86130 0 86186 800 6 wbs_dat_o[18]
port 357 nsew signal output
rlabel metal2 s 89994 0 90050 800 6 wbs_dat_o[19]
port 358 nsew signal output
rlabel metal2 s 16118 0 16174 800 6 wbs_dat_o[1]
port 359 nsew signal output
rlabel metal2 s 93858 0 93914 800 6 wbs_dat_o[20]
port 360 nsew signal output
rlabel metal2 s 97722 0 97778 800 6 wbs_dat_o[21]
port 361 nsew signal output
rlabel metal2 s 101678 0 101734 800 6 wbs_dat_o[22]
port 362 nsew signal output
rlabel metal2 s 105542 0 105598 800 6 wbs_dat_o[23]
port 363 nsew signal output
rlabel metal2 s 109406 0 109462 800 6 wbs_dat_o[24]
port 364 nsew signal output
rlabel metal2 s 113270 0 113326 800 6 wbs_dat_o[25]
port 365 nsew signal output
rlabel metal2 s 117226 0 117282 800 6 wbs_dat_o[26]
port 366 nsew signal output
rlabel metal2 s 121090 0 121146 800 6 wbs_dat_o[27]
port 367 nsew signal output
rlabel metal2 s 124954 0 125010 800 6 wbs_dat_o[28]
port 368 nsew signal output
rlabel metal2 s 128818 0 128874 800 6 wbs_dat_o[29]
port 369 nsew signal output
rlabel metal2 s 21362 0 21418 800 6 wbs_dat_o[2]
port 370 nsew signal output
rlabel metal2 s 132774 0 132830 800 6 wbs_dat_o[30]
port 371 nsew signal output
rlabel metal2 s 136638 0 136694 800 6 wbs_dat_o[31]
port 372 nsew signal output
rlabel metal2 s 26514 0 26570 800 6 wbs_dat_o[3]
port 373 nsew signal output
rlabel metal2 s 31666 0 31722 800 6 wbs_dat_o[4]
port 374 nsew signal output
rlabel metal2 s 35622 0 35678 800 6 wbs_dat_o[5]
port 375 nsew signal output
rlabel metal2 s 39486 0 39542 800 6 wbs_dat_o[6]
port 376 nsew signal output
rlabel metal2 s 43350 0 43406 800 6 wbs_dat_o[7]
port 377 nsew signal output
rlabel metal2 s 47214 0 47270 800 6 wbs_dat_o[8]
port 378 nsew signal output
rlabel metal2 s 51170 0 51226 800 6 wbs_dat_o[9]
port 379 nsew signal output
rlabel metal2 s 12254 0 12310 800 6 wbs_sel_i[0]
port 380 nsew signal input
rlabel metal2 s 17498 0 17554 800 6 wbs_sel_i[1]
port 381 nsew signal input
rlabel metal2 s 22650 0 22706 800 6 wbs_sel_i[2]
port 382 nsew signal input
rlabel metal2 s 27802 0 27858 800 6 wbs_sel_i[3]
port 383 nsew signal input
rlabel metal2 s 5814 0 5870 800 6 wbs_stb_i
port 384 nsew signal input
rlabel metal2 s 7102 0 7158 800 6 wbs_we_i
port 385 nsew signal input
<< properties >>
string LEFclass BLOCK
string FIXED_BBOX 0 0 198125 200269
string LEFview TRUE
string GDS_FILE /local/home/roman/projects/opencircuitdesign/shuttle5/caravel_mpw/openlane/user_proj/runs/user_proj/results/magic/user_proj.gds
string GDS_END 96871328
string GDS_START 1461086
<< end >>

