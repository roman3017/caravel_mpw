magic
tech sky130A
magscale 1 2
timestamp 1643962656
<< obsli1 >>
rect 1104 1445 197679 198033
<< obsm1 >>
rect 1026 620 197691 198756
<< metal2 >>
rect 662 199504 718 200304
rect 1950 199504 2006 200304
rect 3238 199504 3294 200304
rect 4618 199504 4674 200304
rect 5906 199504 5962 200304
rect 7286 199504 7342 200304
rect 8574 199504 8630 200304
rect 9954 199504 10010 200304
rect 11242 199504 11298 200304
rect 12622 199504 12678 200304
rect 13910 199504 13966 200304
rect 15290 199504 15346 200304
rect 16578 199504 16634 200304
rect 17866 199504 17922 200304
rect 19246 199504 19302 200304
rect 20534 199504 20590 200304
rect 21914 199504 21970 200304
rect 23202 199504 23258 200304
rect 24582 199504 24638 200304
rect 25870 199504 25926 200304
rect 27250 199504 27306 200304
rect 28538 199504 28594 200304
rect 29918 199504 29974 200304
rect 31206 199504 31262 200304
rect 32494 199504 32550 200304
rect 33874 199504 33930 200304
rect 35162 199504 35218 200304
rect 36542 199504 36598 200304
rect 37830 199504 37886 200304
rect 39210 199504 39266 200304
rect 40498 199504 40554 200304
rect 41878 199504 41934 200304
rect 43166 199504 43222 200304
rect 44546 199504 44602 200304
rect 45834 199504 45890 200304
rect 47122 199504 47178 200304
rect 48502 199504 48558 200304
rect 49790 199504 49846 200304
rect 51170 199504 51226 200304
rect 52458 199504 52514 200304
rect 53838 199504 53894 200304
rect 55126 199504 55182 200304
rect 56506 199504 56562 200304
rect 57794 199504 57850 200304
rect 59174 199504 59230 200304
rect 60462 199504 60518 200304
rect 61750 199504 61806 200304
rect 63130 199504 63186 200304
rect 64418 199504 64474 200304
rect 65798 199504 65854 200304
rect 67086 199504 67142 200304
rect 68466 199504 68522 200304
rect 69754 199504 69810 200304
rect 71134 199504 71190 200304
rect 72422 199504 72478 200304
rect 73802 199504 73858 200304
rect 75090 199504 75146 200304
rect 76470 199504 76526 200304
rect 77758 199504 77814 200304
rect 79046 199504 79102 200304
rect 80426 199504 80482 200304
rect 81714 199504 81770 200304
rect 83094 199504 83150 200304
rect 84382 199504 84438 200304
rect 85762 199504 85818 200304
rect 87050 199504 87106 200304
rect 88430 199504 88486 200304
rect 89718 199504 89774 200304
rect 91098 199504 91154 200304
rect 92386 199504 92442 200304
rect 93674 199504 93730 200304
rect 95054 199504 95110 200304
rect 96342 199504 96398 200304
rect 97722 199504 97778 200304
rect 99010 199504 99066 200304
rect 100390 199504 100446 200304
rect 101678 199504 101734 200304
rect 103058 199504 103114 200304
rect 104346 199504 104402 200304
rect 105726 199504 105782 200304
rect 107014 199504 107070 200304
rect 108302 199504 108358 200304
rect 109682 199504 109738 200304
rect 110970 199504 111026 200304
rect 112350 199504 112406 200304
rect 113638 199504 113694 200304
rect 115018 199504 115074 200304
rect 116306 199504 116362 200304
rect 117686 199504 117742 200304
rect 118974 199504 119030 200304
rect 120354 199504 120410 200304
rect 121642 199504 121698 200304
rect 122930 199504 122986 200304
rect 124310 199504 124366 200304
rect 125598 199504 125654 200304
rect 126978 199504 127034 200304
rect 128266 199504 128322 200304
rect 129646 199504 129702 200304
rect 130934 199504 130990 200304
rect 132314 199504 132370 200304
rect 133602 199504 133658 200304
rect 134982 199504 135038 200304
rect 136270 199504 136326 200304
rect 137650 199504 137706 200304
rect 138938 199504 138994 200304
rect 140226 199504 140282 200304
rect 141606 199504 141662 200304
rect 142894 199504 142950 200304
rect 144274 199504 144330 200304
rect 145562 199504 145618 200304
rect 146942 199504 146998 200304
rect 148230 199504 148286 200304
rect 149610 199504 149666 200304
rect 150898 199504 150954 200304
rect 152278 199504 152334 200304
rect 153566 199504 153622 200304
rect 154854 199504 154910 200304
rect 156234 199504 156290 200304
rect 157522 199504 157578 200304
rect 158902 199504 158958 200304
rect 160190 199504 160246 200304
rect 161570 199504 161626 200304
rect 162858 199504 162914 200304
rect 164238 199504 164294 200304
rect 165526 199504 165582 200304
rect 166906 199504 166962 200304
rect 168194 199504 168250 200304
rect 169482 199504 169538 200304
rect 170862 199504 170918 200304
rect 172150 199504 172206 200304
rect 173530 199504 173586 200304
rect 174818 199504 174874 200304
rect 176198 199504 176254 200304
rect 177486 199504 177542 200304
rect 178866 199504 178922 200304
rect 180154 199504 180210 200304
rect 181534 199504 181590 200304
rect 182822 199504 182878 200304
rect 184110 199504 184166 200304
rect 185490 199504 185546 200304
rect 186778 199504 186834 200304
rect 188158 199504 188214 200304
rect 189446 199504 189502 200304
rect 190826 199504 190882 200304
rect 192114 199504 192170 200304
rect 193494 199504 193550 200304
rect 194782 199504 194838 200304
rect 196162 199504 196218 200304
rect 197450 199504 197506 200304
rect 570 0 626 800
rect 1766 0 1822 800
rect 3054 0 3110 800
rect 4342 0 4398 800
rect 5630 0 5686 800
rect 6918 0 6974 800
rect 8206 0 8262 800
rect 9494 0 9550 800
rect 10782 0 10838 800
rect 12070 0 12126 800
rect 13266 0 13322 800
rect 14554 0 14610 800
rect 15842 0 15898 800
rect 17130 0 17186 800
rect 18418 0 18474 800
rect 19706 0 19762 800
rect 20994 0 21050 800
rect 22282 0 22338 800
rect 23570 0 23626 800
rect 24858 0 24914 800
rect 26054 0 26110 800
rect 27342 0 27398 800
rect 28630 0 28686 800
rect 29918 0 29974 800
rect 31206 0 31262 800
rect 32494 0 32550 800
rect 33782 0 33838 800
rect 35070 0 35126 800
rect 36358 0 36414 800
rect 37646 0 37702 800
rect 38842 0 38898 800
rect 40130 0 40186 800
rect 41418 0 41474 800
rect 42706 0 42762 800
rect 43994 0 44050 800
rect 45282 0 45338 800
rect 46570 0 46626 800
rect 47858 0 47914 800
rect 49146 0 49202 800
rect 50342 0 50398 800
rect 51630 0 51686 800
rect 52918 0 52974 800
rect 54206 0 54262 800
rect 55494 0 55550 800
rect 56782 0 56838 800
rect 58070 0 58126 800
rect 59358 0 59414 800
rect 60646 0 60702 800
rect 61934 0 61990 800
rect 63130 0 63186 800
rect 64418 0 64474 800
rect 65706 0 65762 800
rect 66994 0 67050 800
rect 68282 0 68338 800
rect 69570 0 69626 800
rect 70858 0 70914 800
rect 72146 0 72202 800
rect 73434 0 73490 800
rect 74722 0 74778 800
rect 75918 0 75974 800
rect 77206 0 77262 800
rect 78494 0 78550 800
rect 79782 0 79838 800
rect 81070 0 81126 800
rect 82358 0 82414 800
rect 83646 0 83702 800
rect 84934 0 84990 800
rect 86222 0 86278 800
rect 87418 0 87474 800
rect 88706 0 88762 800
rect 89994 0 90050 800
rect 91282 0 91338 800
rect 92570 0 92626 800
rect 93858 0 93914 800
rect 95146 0 95202 800
rect 96434 0 96490 800
rect 97722 0 97778 800
rect 99010 0 99066 800
rect 100206 0 100262 800
rect 101494 0 101550 800
rect 102782 0 102838 800
rect 104070 0 104126 800
rect 105358 0 105414 800
rect 106646 0 106702 800
rect 107934 0 107990 800
rect 109222 0 109278 800
rect 110510 0 110566 800
rect 111798 0 111854 800
rect 112994 0 113050 800
rect 114282 0 114338 800
rect 115570 0 115626 800
rect 116858 0 116914 800
rect 118146 0 118202 800
rect 119434 0 119490 800
rect 120722 0 120778 800
rect 122010 0 122066 800
rect 123298 0 123354 800
rect 124494 0 124550 800
rect 125782 0 125838 800
rect 127070 0 127126 800
rect 128358 0 128414 800
rect 129646 0 129702 800
rect 130934 0 130990 800
rect 132222 0 132278 800
rect 133510 0 133566 800
rect 134798 0 134854 800
rect 136086 0 136142 800
rect 137282 0 137338 800
rect 138570 0 138626 800
rect 139858 0 139914 800
rect 141146 0 141202 800
rect 142434 0 142490 800
rect 143722 0 143778 800
rect 145010 0 145066 800
rect 146298 0 146354 800
rect 147586 0 147642 800
rect 148874 0 148930 800
rect 150070 0 150126 800
rect 151358 0 151414 800
rect 152646 0 152702 800
rect 153934 0 153990 800
rect 155222 0 155278 800
rect 156510 0 156566 800
rect 157798 0 157854 800
rect 159086 0 159142 800
rect 160374 0 160430 800
rect 161570 0 161626 800
rect 162858 0 162914 800
rect 164146 0 164202 800
rect 165434 0 165490 800
rect 166722 0 166778 800
rect 168010 0 168066 800
rect 169298 0 169354 800
rect 170586 0 170642 800
rect 171874 0 171930 800
rect 173162 0 173218 800
rect 174358 0 174414 800
rect 175646 0 175702 800
rect 176934 0 176990 800
rect 178222 0 178278 800
rect 179510 0 179566 800
rect 180798 0 180854 800
rect 182086 0 182142 800
rect 183374 0 183430 800
rect 184662 0 184718 800
rect 185950 0 186006 800
rect 187146 0 187202 800
rect 188434 0 188490 800
rect 189722 0 189778 800
rect 191010 0 191066 800
rect 192298 0 192354 800
rect 193586 0 193642 800
rect 194874 0 194930 800
rect 196162 0 196218 800
rect 197450 0 197506 800
<< obsm2 >>
rect 110 199448 606 199594
rect 774 199448 1894 199594
rect 2062 199448 3182 199594
rect 3350 199448 4562 199594
rect 4730 199448 5850 199594
rect 6018 199448 7230 199594
rect 7398 199448 8518 199594
rect 8686 199448 9898 199594
rect 10066 199448 11186 199594
rect 11354 199448 12566 199594
rect 12734 199448 13854 199594
rect 14022 199448 15234 199594
rect 15402 199448 16522 199594
rect 16690 199448 17810 199594
rect 17978 199448 19190 199594
rect 19358 199448 20478 199594
rect 20646 199448 21858 199594
rect 22026 199448 23146 199594
rect 23314 199448 24526 199594
rect 24694 199448 25814 199594
rect 25982 199448 27194 199594
rect 27362 199448 28482 199594
rect 28650 199448 29862 199594
rect 30030 199448 31150 199594
rect 31318 199448 32438 199594
rect 32606 199448 33818 199594
rect 33986 199448 35106 199594
rect 35274 199448 36486 199594
rect 36654 199448 37774 199594
rect 37942 199448 39154 199594
rect 39322 199448 40442 199594
rect 40610 199448 41822 199594
rect 41990 199448 43110 199594
rect 43278 199448 44490 199594
rect 44658 199448 45778 199594
rect 45946 199448 47066 199594
rect 47234 199448 48446 199594
rect 48614 199448 49734 199594
rect 49902 199448 51114 199594
rect 51282 199448 52402 199594
rect 52570 199448 53782 199594
rect 53950 199448 55070 199594
rect 55238 199448 56450 199594
rect 56618 199448 57738 199594
rect 57906 199448 59118 199594
rect 59286 199448 60406 199594
rect 60574 199448 61694 199594
rect 61862 199448 63074 199594
rect 63242 199448 64362 199594
rect 64530 199448 65742 199594
rect 65910 199448 67030 199594
rect 67198 199448 68410 199594
rect 68578 199448 69698 199594
rect 69866 199448 71078 199594
rect 71246 199448 72366 199594
rect 72534 199448 73746 199594
rect 73914 199448 75034 199594
rect 75202 199448 76414 199594
rect 76582 199448 77702 199594
rect 77870 199448 78990 199594
rect 79158 199448 80370 199594
rect 80538 199448 81658 199594
rect 81826 199448 83038 199594
rect 83206 199448 84326 199594
rect 84494 199448 85706 199594
rect 85874 199448 86994 199594
rect 87162 199448 88374 199594
rect 88542 199448 89662 199594
rect 89830 199448 91042 199594
rect 91210 199448 92330 199594
rect 92498 199448 93618 199594
rect 93786 199448 94998 199594
rect 95166 199448 96286 199594
rect 96454 199448 97666 199594
rect 97834 199448 98954 199594
rect 99122 199448 100334 199594
rect 100502 199448 101622 199594
rect 101790 199448 103002 199594
rect 103170 199448 104290 199594
rect 104458 199448 105670 199594
rect 105838 199448 106958 199594
rect 107126 199448 108246 199594
rect 108414 199448 109626 199594
rect 109794 199448 110914 199594
rect 111082 199448 112294 199594
rect 112462 199448 113582 199594
rect 113750 199448 114962 199594
rect 115130 199448 116250 199594
rect 116418 199448 117630 199594
rect 117798 199448 118918 199594
rect 119086 199448 120298 199594
rect 120466 199448 121586 199594
rect 121754 199448 122874 199594
rect 123042 199448 124254 199594
rect 124422 199448 125542 199594
rect 125710 199448 126922 199594
rect 127090 199448 128210 199594
rect 128378 199448 129590 199594
rect 129758 199448 130878 199594
rect 131046 199448 132258 199594
rect 132426 199448 133546 199594
rect 133714 199448 134926 199594
rect 135094 199448 136214 199594
rect 136382 199448 137594 199594
rect 137762 199448 138882 199594
rect 139050 199448 140170 199594
rect 140338 199448 141550 199594
rect 141718 199448 142838 199594
rect 143006 199448 144218 199594
rect 144386 199448 145506 199594
rect 145674 199448 146886 199594
rect 147054 199448 148174 199594
rect 148342 199448 149554 199594
rect 149722 199448 150842 199594
rect 151010 199448 152222 199594
rect 152390 199448 153510 199594
rect 153678 199448 154798 199594
rect 154966 199448 156178 199594
rect 156346 199448 157466 199594
rect 157634 199448 158846 199594
rect 159014 199448 160134 199594
rect 160302 199448 161514 199594
rect 161682 199448 162802 199594
rect 162970 199448 164182 199594
rect 164350 199448 165470 199594
rect 165638 199448 166850 199594
rect 167018 199448 168138 199594
rect 168306 199448 169426 199594
rect 169594 199448 170806 199594
rect 170974 199448 172094 199594
rect 172262 199448 173474 199594
rect 173642 199448 174762 199594
rect 174930 199448 176142 199594
rect 176310 199448 177430 199594
rect 177598 199448 178810 199594
rect 178978 199448 180098 199594
rect 180266 199448 181478 199594
rect 181646 199448 182766 199594
rect 182934 199448 184054 199594
rect 184222 199448 185434 199594
rect 185602 199448 186722 199594
rect 186890 199448 188102 199594
rect 188270 199448 189390 199594
rect 189558 199448 190770 199594
rect 190938 199448 192058 199594
rect 192226 199448 193438 199594
rect 193606 199448 194726 199594
rect 194894 199448 196106 199594
rect 196274 199448 197394 199594
rect 110 856 197504 199448
rect 110 614 514 856
rect 682 614 1710 856
rect 1878 614 2998 856
rect 3166 614 4286 856
rect 4454 614 5574 856
rect 5742 614 6862 856
rect 7030 614 8150 856
rect 8318 614 9438 856
rect 9606 614 10726 856
rect 10894 614 12014 856
rect 12182 614 13210 856
rect 13378 614 14498 856
rect 14666 614 15786 856
rect 15954 614 17074 856
rect 17242 614 18362 856
rect 18530 614 19650 856
rect 19818 614 20938 856
rect 21106 614 22226 856
rect 22394 614 23514 856
rect 23682 614 24802 856
rect 24970 614 25998 856
rect 26166 614 27286 856
rect 27454 614 28574 856
rect 28742 614 29862 856
rect 30030 614 31150 856
rect 31318 614 32438 856
rect 32606 614 33726 856
rect 33894 614 35014 856
rect 35182 614 36302 856
rect 36470 614 37590 856
rect 37758 614 38786 856
rect 38954 614 40074 856
rect 40242 614 41362 856
rect 41530 614 42650 856
rect 42818 614 43938 856
rect 44106 614 45226 856
rect 45394 614 46514 856
rect 46682 614 47802 856
rect 47970 614 49090 856
rect 49258 614 50286 856
rect 50454 614 51574 856
rect 51742 614 52862 856
rect 53030 614 54150 856
rect 54318 614 55438 856
rect 55606 614 56726 856
rect 56894 614 58014 856
rect 58182 614 59302 856
rect 59470 614 60590 856
rect 60758 614 61878 856
rect 62046 614 63074 856
rect 63242 614 64362 856
rect 64530 614 65650 856
rect 65818 614 66938 856
rect 67106 614 68226 856
rect 68394 614 69514 856
rect 69682 614 70802 856
rect 70970 614 72090 856
rect 72258 614 73378 856
rect 73546 614 74666 856
rect 74834 614 75862 856
rect 76030 614 77150 856
rect 77318 614 78438 856
rect 78606 614 79726 856
rect 79894 614 81014 856
rect 81182 614 82302 856
rect 82470 614 83590 856
rect 83758 614 84878 856
rect 85046 614 86166 856
rect 86334 614 87362 856
rect 87530 614 88650 856
rect 88818 614 89938 856
rect 90106 614 91226 856
rect 91394 614 92514 856
rect 92682 614 93802 856
rect 93970 614 95090 856
rect 95258 614 96378 856
rect 96546 614 97666 856
rect 97834 614 98954 856
rect 99122 614 100150 856
rect 100318 614 101438 856
rect 101606 614 102726 856
rect 102894 614 104014 856
rect 104182 614 105302 856
rect 105470 614 106590 856
rect 106758 614 107878 856
rect 108046 614 109166 856
rect 109334 614 110454 856
rect 110622 614 111742 856
rect 111910 614 112938 856
rect 113106 614 114226 856
rect 114394 614 115514 856
rect 115682 614 116802 856
rect 116970 614 118090 856
rect 118258 614 119378 856
rect 119546 614 120666 856
rect 120834 614 121954 856
rect 122122 614 123242 856
rect 123410 614 124438 856
rect 124606 614 125726 856
rect 125894 614 127014 856
rect 127182 614 128302 856
rect 128470 614 129590 856
rect 129758 614 130878 856
rect 131046 614 132166 856
rect 132334 614 133454 856
rect 133622 614 134742 856
rect 134910 614 136030 856
rect 136198 614 137226 856
rect 137394 614 138514 856
rect 138682 614 139802 856
rect 139970 614 141090 856
rect 141258 614 142378 856
rect 142546 614 143666 856
rect 143834 614 144954 856
rect 145122 614 146242 856
rect 146410 614 147530 856
rect 147698 614 148818 856
rect 148986 614 150014 856
rect 150182 614 151302 856
rect 151470 614 152590 856
rect 152758 614 153878 856
rect 154046 614 155166 856
rect 155334 614 156454 856
rect 156622 614 157742 856
rect 157910 614 159030 856
rect 159198 614 160318 856
rect 160486 614 161514 856
rect 161682 614 162802 856
rect 162970 614 164090 856
rect 164258 614 165378 856
rect 165546 614 166666 856
rect 166834 614 167954 856
rect 168122 614 169242 856
rect 169410 614 170530 856
rect 170698 614 171818 856
rect 171986 614 173106 856
rect 173274 614 174302 856
rect 174470 614 175590 856
rect 175758 614 176878 856
rect 177046 614 178166 856
rect 178334 614 179454 856
rect 179622 614 180742 856
rect 180910 614 182030 856
rect 182198 614 183318 856
rect 183486 614 184606 856
rect 184774 614 185894 856
rect 186062 614 187090 856
rect 187258 614 188378 856
rect 188546 614 189666 856
rect 189834 614 190954 856
rect 191122 614 192242 856
rect 192410 614 193530 856
rect 193698 614 194818 856
rect 194986 614 196106 856
rect 196274 614 197394 856
<< metal3 >>
rect 0 197752 800 197872
rect 197360 197480 198160 197600
rect 0 192992 800 193112
rect 197360 192040 198160 192160
rect 0 188232 800 188352
rect 197360 186600 198160 186720
rect 0 183472 800 183592
rect 197360 181160 198160 181280
rect 0 178712 800 178832
rect 197360 175720 198160 175840
rect 0 173952 800 174072
rect 197360 170416 198160 170536
rect 0 169192 800 169312
rect 197360 164976 198160 165096
rect 0 164432 800 164552
rect 0 159672 800 159792
rect 197360 159536 198160 159656
rect 0 154912 800 155032
rect 197360 154096 198160 154216
rect 0 150152 800 150272
rect 197360 148656 198160 148776
rect 0 145392 800 145512
rect 197360 143352 198160 143472
rect 0 140632 800 140752
rect 197360 137912 198160 138032
rect 0 135872 800 135992
rect 197360 132472 198160 132592
rect 0 130976 800 131096
rect 197360 127032 198160 127152
rect 0 126216 800 126336
rect 0 121456 800 121576
rect 197360 121592 198160 121712
rect 0 116696 800 116816
rect 197360 116288 198160 116408
rect 0 111936 800 112056
rect 197360 110848 198160 110968
rect 0 107176 800 107296
rect 197360 105408 198160 105528
rect 0 102416 800 102536
rect 197360 99968 198160 100088
rect 0 97656 800 97776
rect 197360 94528 198160 94648
rect 0 92896 800 93016
rect 197360 89088 198160 89208
rect 0 88136 800 88256
rect 197360 83784 198160 83904
rect 0 83376 800 83496
rect 0 78616 800 78736
rect 197360 78344 198160 78464
rect 0 73856 800 73976
rect 197360 72904 198160 73024
rect 0 69096 800 69216
rect 197360 67464 198160 67584
rect 0 64200 800 64320
rect 197360 62024 198160 62144
rect 0 59440 800 59560
rect 197360 56720 198160 56840
rect 0 54680 800 54800
rect 197360 51280 198160 51400
rect 0 49920 800 50040
rect 197360 45840 198160 45960
rect 0 45160 800 45280
rect 0 40400 800 40520
rect 197360 40400 198160 40520
rect 0 35640 800 35760
rect 197360 34960 198160 35080
rect 0 30880 800 31000
rect 197360 29656 198160 29776
rect 0 26120 800 26240
rect 197360 24216 198160 24336
rect 0 21360 800 21480
rect 197360 18776 198160 18896
rect 0 16600 800 16720
rect 197360 13336 198160 13456
rect 0 11840 800 11960
rect 197360 7896 198160 8016
rect 0 7080 800 7200
rect 197360 2592 198160 2712
rect 0 2320 800 2440
<< obsm3 >>
rect 105 197952 197360 198253
rect 880 197680 197360 197952
rect 880 197672 197280 197680
rect 105 197400 197280 197672
rect 105 193192 197360 197400
rect 880 192912 197360 193192
rect 105 192240 197360 192912
rect 105 191960 197280 192240
rect 105 188432 197360 191960
rect 880 188152 197360 188432
rect 105 186800 197360 188152
rect 105 186520 197280 186800
rect 105 183672 197360 186520
rect 880 183392 197360 183672
rect 105 181360 197360 183392
rect 105 181080 197280 181360
rect 105 178912 197360 181080
rect 880 178632 197360 178912
rect 105 175920 197360 178632
rect 105 175640 197280 175920
rect 105 174152 197360 175640
rect 880 173872 197360 174152
rect 105 170616 197360 173872
rect 105 170336 197280 170616
rect 105 169392 197360 170336
rect 880 169112 197360 169392
rect 105 165176 197360 169112
rect 105 164896 197280 165176
rect 105 164632 197360 164896
rect 880 164352 197360 164632
rect 105 159872 197360 164352
rect 880 159736 197360 159872
rect 880 159592 197280 159736
rect 105 159456 197280 159592
rect 105 155112 197360 159456
rect 880 154832 197360 155112
rect 105 154296 197360 154832
rect 105 154016 197280 154296
rect 105 150352 197360 154016
rect 880 150072 197360 150352
rect 105 148856 197360 150072
rect 105 148576 197280 148856
rect 105 145592 197360 148576
rect 880 145312 197360 145592
rect 105 143552 197360 145312
rect 105 143272 197280 143552
rect 105 140832 197360 143272
rect 880 140552 197360 140832
rect 105 138112 197360 140552
rect 105 137832 197280 138112
rect 105 136072 197360 137832
rect 880 135792 197360 136072
rect 105 132672 197360 135792
rect 105 132392 197280 132672
rect 105 131176 197360 132392
rect 880 130896 197360 131176
rect 105 127232 197360 130896
rect 105 126952 197280 127232
rect 105 126416 197360 126952
rect 880 126136 197360 126416
rect 105 121792 197360 126136
rect 105 121656 197280 121792
rect 880 121512 197280 121656
rect 880 121376 197360 121512
rect 105 116896 197360 121376
rect 880 116616 197360 116896
rect 105 116488 197360 116616
rect 105 116208 197280 116488
rect 105 112136 197360 116208
rect 880 111856 197360 112136
rect 105 111048 197360 111856
rect 105 110768 197280 111048
rect 105 107376 197360 110768
rect 880 107096 197360 107376
rect 105 105608 197360 107096
rect 105 105328 197280 105608
rect 105 102616 197360 105328
rect 880 102336 197360 102616
rect 105 100168 197360 102336
rect 105 99888 197280 100168
rect 105 97856 197360 99888
rect 880 97576 197360 97856
rect 105 94728 197360 97576
rect 105 94448 197280 94728
rect 105 93096 197360 94448
rect 880 92816 197360 93096
rect 105 89288 197360 92816
rect 105 89008 197280 89288
rect 105 88336 197360 89008
rect 880 88056 197360 88336
rect 105 83984 197360 88056
rect 105 83704 197280 83984
rect 105 83576 197360 83704
rect 880 83296 197360 83576
rect 105 78816 197360 83296
rect 880 78544 197360 78816
rect 880 78536 197280 78544
rect 105 78264 197280 78536
rect 105 74056 197360 78264
rect 880 73776 197360 74056
rect 105 73104 197360 73776
rect 105 72824 197280 73104
rect 105 69296 197360 72824
rect 880 69016 197360 69296
rect 105 67664 197360 69016
rect 105 67384 197280 67664
rect 105 64400 197360 67384
rect 880 64120 197360 64400
rect 105 62224 197360 64120
rect 105 61944 197280 62224
rect 105 59640 197360 61944
rect 880 59360 197360 59640
rect 105 56920 197360 59360
rect 105 56640 197280 56920
rect 105 54880 197360 56640
rect 880 54600 197360 54880
rect 105 51480 197360 54600
rect 105 51200 197280 51480
rect 105 50120 197360 51200
rect 880 49840 197360 50120
rect 105 46040 197360 49840
rect 105 45760 197280 46040
rect 105 45360 197360 45760
rect 880 45080 197360 45360
rect 105 40600 197360 45080
rect 880 40320 197280 40600
rect 105 35840 197360 40320
rect 880 35560 197360 35840
rect 105 35160 197360 35560
rect 105 34880 197280 35160
rect 105 31080 197360 34880
rect 880 30800 197360 31080
rect 105 29856 197360 30800
rect 105 29576 197280 29856
rect 105 26320 197360 29576
rect 880 26040 197360 26320
rect 105 24416 197360 26040
rect 105 24136 197280 24416
rect 105 21560 197360 24136
rect 880 21280 197360 21560
rect 105 18976 197360 21280
rect 105 18696 197280 18976
rect 105 16800 197360 18696
rect 880 16520 197360 16800
rect 105 13536 197360 16520
rect 105 13256 197280 13536
rect 105 12040 197360 13256
rect 880 11760 197360 12040
rect 105 8096 197360 11760
rect 105 7816 197280 8096
rect 105 7280 197360 7816
rect 880 7000 197360 7280
rect 105 2792 197360 7000
rect 105 2520 197280 2792
rect 880 2512 197280 2520
rect 880 2240 197360 2512
rect 105 1803 197360 2240
<< metal4 >>
rect 4208 2128 4528 198064
rect 19568 2128 19888 198064
rect 34928 2128 35248 198064
rect 50288 2128 50608 198064
rect 65648 2128 65968 198064
rect 81008 2128 81328 198064
rect 96368 2128 96688 198064
rect 111728 2128 112048 198064
rect 127088 2128 127408 198064
rect 142448 2128 142768 198064
rect 157808 2128 158128 198064
rect 173168 2128 173488 198064
rect 188528 2128 188848 198064
<< obsm4 >>
rect 40539 198144 195533 198253
rect 40539 5883 50208 198144
rect 50688 5883 65568 198144
rect 66048 5883 80928 198144
rect 81408 5883 96288 198144
rect 96768 5883 111648 198144
rect 112128 5883 127008 198144
rect 127488 5883 142368 198144
rect 142848 5883 157728 198144
rect 158208 5883 173088 198144
rect 173568 5883 188448 198144
rect 188928 5883 195533 198144
<< labels >>
rlabel metal3 s 0 2320 800 2440 6 clk_i
port 1 nsew signal input
rlabel metal3 s 0 11840 800 11960 6 i_dout0[0]
port 2 nsew signal input
rlabel metal2 s 170862 199504 170918 200304 6 i_dout0[10]
port 3 nsew signal input
rlabel metal3 s 0 92896 800 93016 6 i_dout0[11]
port 4 nsew signal input
rlabel metal3 s 197360 116288 198160 116408 6 i_dout0[12]
port 5 nsew signal input
rlabel metal2 s 172150 199504 172206 200304 6 i_dout0[13]
port 6 nsew signal input
rlabel metal3 s 0 121456 800 121576 6 i_dout0[14]
port 7 nsew signal input
rlabel metal3 s 0 126216 800 126336 6 i_dout0[15]
port 8 nsew signal input
rlabel metal2 s 176198 199504 176254 200304 6 i_dout0[16]
port 9 nsew signal input
rlabel metal3 s 197360 137912 198160 138032 6 i_dout0[17]
port 10 nsew signal input
rlabel metal3 s 0 140632 800 140752 6 i_dout0[18]
port 11 nsew signal input
rlabel metal3 s 0 150152 800 150272 6 i_dout0[19]
port 12 nsew signal input
rlabel metal3 s 0 16600 800 16720 6 i_dout0[1]
port 13 nsew signal input
rlabel metal3 s 0 159672 800 159792 6 i_dout0[20]
port 14 nsew signal input
rlabel metal2 s 181534 199504 181590 200304 6 i_dout0[21]
port 15 nsew signal input
rlabel metal2 s 180798 0 180854 800 6 i_dout0[22]
port 16 nsew signal input
rlabel metal3 s 197360 159536 198160 159656 6 i_dout0[23]
port 17 nsew signal input
rlabel metal2 s 182086 0 182142 800 6 i_dout0[24]
port 18 nsew signal input
rlabel metal3 s 0 178712 800 178832 6 i_dout0[25]
port 19 nsew signal input
rlabel metal2 s 188434 0 188490 800 6 i_dout0[26]
port 20 nsew signal input
rlabel metal2 s 191010 0 191066 800 6 i_dout0[27]
port 21 nsew signal input
rlabel metal3 s 197360 181160 198160 181280 6 i_dout0[28]
port 22 nsew signal input
rlabel metal3 s 0 197752 800 197872 6 i_dout0[29]
port 23 nsew signal input
rlabel metal2 s 156234 199504 156290 200304 6 i_dout0[2]
port 24 nsew signal input
rlabel metal2 s 193494 199504 193550 200304 6 i_dout0[30]
port 25 nsew signal input
rlabel metal2 s 197450 0 197506 800 6 i_dout0[31]
port 26 nsew signal input
rlabel metal3 s 197360 62024 198160 62144 6 i_dout0[3]
port 27 nsew signal input
rlabel metal2 s 152646 0 152702 800 6 i_dout0[4]
port 28 nsew signal input
rlabel metal3 s 0 59440 800 59560 6 i_dout0[5]
port 29 nsew signal input
rlabel metal2 s 159086 0 159142 800 6 i_dout0[6]
port 30 nsew signal input
rlabel metal3 s 197360 89088 198160 89208 6 i_dout0[7]
port 31 nsew signal input
rlabel metal2 s 164146 0 164202 800 6 i_dout0[8]
port 32 nsew signal input
rlabel metal2 s 165526 199504 165582 200304 6 i_dout0[9]
port 33 nsew signal input
rlabel metal2 s 152278 199504 152334 200304 6 i_dout0_1[0]
port 34 nsew signal input
rlabel metal2 s 169482 199504 169538 200304 6 i_dout0_1[10]
port 35 nsew signal input
rlabel metal3 s 0 88136 800 88256 6 i_dout0_1[11]
port 36 nsew signal input
rlabel metal3 s 0 102416 800 102536 6 i_dout0_1[12]
port 37 nsew signal input
rlabel metal3 s 0 107176 800 107296 6 i_dout0_1[13]
port 38 nsew signal input
rlabel metal2 s 171874 0 171930 800 6 i_dout0_1[14]
port 39 nsew signal input
rlabel metal2 s 174818 199504 174874 200304 6 i_dout0_1[15]
port 40 nsew signal input
rlabel metal3 s 197360 127032 198160 127152 6 i_dout0_1[16]
port 41 nsew signal input
rlabel metal2 s 177486 199504 177542 200304 6 i_dout0_1[17]
port 42 nsew signal input
rlabel metal3 s 0 135872 800 135992 6 i_dout0_1[18]
port 43 nsew signal input
rlabel metal2 s 178866 199504 178922 200304 6 i_dout0_1[19]
port 44 nsew signal input
rlabel metal3 s 197360 29656 198160 29776 6 i_dout0_1[1]
port 45 nsew signal input
rlabel metal3 s 0 154912 800 155032 6 i_dout0_1[20]
port 46 nsew signal input
rlabel metal2 s 179510 0 179566 800 6 i_dout0_1[21]
port 47 nsew signal input
rlabel metal2 s 184110 199504 184166 200304 6 i_dout0_1[22]
port 48 nsew signal input
rlabel metal2 s 186778 199504 186834 200304 6 i_dout0_1[23]
port 49 nsew signal input
rlabel metal2 s 188158 199504 188214 200304 6 i_dout0_1[24]
port 50 nsew signal input
rlabel metal2 s 189446 199504 189502 200304 6 i_dout0_1[25]
port 51 nsew signal input
rlabel metal3 s 197360 170416 198160 170536 6 i_dout0_1[26]
port 52 nsew signal input
rlabel metal3 s 197360 175720 198160 175840 6 i_dout0_1[27]
port 53 nsew signal input
rlabel metal2 s 193586 0 193642 800 6 i_dout0_1[28]
port 54 nsew signal input
rlabel metal3 s 0 192992 800 193112 6 i_dout0_1[29]
port 55 nsew signal input
rlabel metal3 s 0 26120 800 26240 6 i_dout0_1[2]
port 56 nsew signal input
rlabel metal3 s 197360 192040 198160 192160 6 i_dout0_1[30]
port 57 nsew signal input
rlabel metal3 s 197360 197480 198160 197600 6 i_dout0_1[31]
port 58 nsew signal input
rlabel metal3 s 197360 56720 198160 56840 6 i_dout0_1[3]
port 59 nsew signal input
rlabel metal3 s 0 49920 800 50040 6 i_dout0_1[4]
port 60 nsew signal input
rlabel metal2 s 158902 199504 158958 200304 6 i_dout0_1[5]
port 61 nsew signal input
rlabel metal2 s 157798 0 157854 800 6 i_dout0_1[6]
port 62 nsew signal input
rlabel metal2 s 162858 0 162914 800 6 i_dout0_1[7]
port 63 nsew signal input
rlabel metal3 s 0 83376 800 83496 6 i_dout0_1[8]
port 64 nsew signal input
rlabel metal2 s 164238 199504 164294 200304 6 i_dout0_1[9]
port 65 nsew signal input
rlabel metal2 s 662 199504 718 200304 6 io_in[0]
port 66 nsew signal input
rlabel metal2 s 40498 199504 40554 200304 6 io_in[10]
port 67 nsew signal input
rlabel metal2 s 44546 199504 44602 200304 6 io_in[11]
port 68 nsew signal input
rlabel metal2 s 48502 199504 48558 200304 6 io_in[12]
port 69 nsew signal input
rlabel metal2 s 52458 199504 52514 200304 6 io_in[13]
port 70 nsew signal input
rlabel metal2 s 56506 199504 56562 200304 6 io_in[14]
port 71 nsew signal input
rlabel metal2 s 60462 199504 60518 200304 6 io_in[15]
port 72 nsew signal input
rlabel metal2 s 64418 199504 64474 200304 6 io_in[16]
port 73 nsew signal input
rlabel metal2 s 68466 199504 68522 200304 6 io_in[17]
port 74 nsew signal input
rlabel metal2 s 72422 199504 72478 200304 6 io_in[18]
port 75 nsew signal input
rlabel metal2 s 76470 199504 76526 200304 6 io_in[19]
port 76 nsew signal input
rlabel metal2 s 4618 199504 4674 200304 6 io_in[1]
port 77 nsew signal input
rlabel metal2 s 80426 199504 80482 200304 6 io_in[20]
port 78 nsew signal input
rlabel metal2 s 84382 199504 84438 200304 6 io_in[21]
port 79 nsew signal input
rlabel metal2 s 88430 199504 88486 200304 6 io_in[22]
port 80 nsew signal input
rlabel metal2 s 92386 199504 92442 200304 6 io_in[23]
port 81 nsew signal input
rlabel metal2 s 96342 199504 96398 200304 6 io_in[24]
port 82 nsew signal input
rlabel metal2 s 100390 199504 100446 200304 6 io_in[25]
port 83 nsew signal input
rlabel metal2 s 104346 199504 104402 200304 6 io_in[26]
port 84 nsew signal input
rlabel metal2 s 108302 199504 108358 200304 6 io_in[27]
port 85 nsew signal input
rlabel metal2 s 112350 199504 112406 200304 6 io_in[28]
port 86 nsew signal input
rlabel metal2 s 116306 199504 116362 200304 6 io_in[29]
port 87 nsew signal input
rlabel metal2 s 8574 199504 8630 200304 6 io_in[2]
port 88 nsew signal input
rlabel metal2 s 120354 199504 120410 200304 6 io_in[30]
port 89 nsew signal input
rlabel metal2 s 124310 199504 124366 200304 6 io_in[31]
port 90 nsew signal input
rlabel metal2 s 128266 199504 128322 200304 6 io_in[32]
port 91 nsew signal input
rlabel metal2 s 132314 199504 132370 200304 6 io_in[33]
port 92 nsew signal input
rlabel metal2 s 136270 199504 136326 200304 6 io_in[34]
port 93 nsew signal input
rlabel metal2 s 140226 199504 140282 200304 6 io_in[35]
port 94 nsew signal input
rlabel metal2 s 144274 199504 144330 200304 6 io_in[36]
port 95 nsew signal input
rlabel metal2 s 148230 199504 148286 200304 6 io_in[37]
port 96 nsew signal input
rlabel metal2 s 12622 199504 12678 200304 6 io_in[3]
port 97 nsew signal input
rlabel metal2 s 16578 199504 16634 200304 6 io_in[4]
port 98 nsew signal input
rlabel metal2 s 20534 199504 20590 200304 6 io_in[5]
port 99 nsew signal input
rlabel metal2 s 24582 199504 24638 200304 6 io_in[6]
port 100 nsew signal input
rlabel metal2 s 28538 199504 28594 200304 6 io_in[7]
port 101 nsew signal input
rlabel metal2 s 32494 199504 32550 200304 6 io_in[8]
port 102 nsew signal input
rlabel metal2 s 36542 199504 36598 200304 6 io_in[9]
port 103 nsew signal input
rlabel metal2 s 1950 199504 2006 200304 6 io_oeb[0]
port 104 nsew signal output
rlabel metal2 s 41878 199504 41934 200304 6 io_oeb[10]
port 105 nsew signal output
rlabel metal2 s 45834 199504 45890 200304 6 io_oeb[11]
port 106 nsew signal output
rlabel metal2 s 49790 199504 49846 200304 6 io_oeb[12]
port 107 nsew signal output
rlabel metal2 s 53838 199504 53894 200304 6 io_oeb[13]
port 108 nsew signal output
rlabel metal2 s 57794 199504 57850 200304 6 io_oeb[14]
port 109 nsew signal output
rlabel metal2 s 61750 199504 61806 200304 6 io_oeb[15]
port 110 nsew signal output
rlabel metal2 s 65798 199504 65854 200304 6 io_oeb[16]
port 111 nsew signal output
rlabel metal2 s 69754 199504 69810 200304 6 io_oeb[17]
port 112 nsew signal output
rlabel metal2 s 73802 199504 73858 200304 6 io_oeb[18]
port 113 nsew signal output
rlabel metal2 s 77758 199504 77814 200304 6 io_oeb[19]
port 114 nsew signal output
rlabel metal2 s 5906 199504 5962 200304 6 io_oeb[1]
port 115 nsew signal output
rlabel metal2 s 81714 199504 81770 200304 6 io_oeb[20]
port 116 nsew signal output
rlabel metal2 s 85762 199504 85818 200304 6 io_oeb[21]
port 117 nsew signal output
rlabel metal2 s 89718 199504 89774 200304 6 io_oeb[22]
port 118 nsew signal output
rlabel metal2 s 93674 199504 93730 200304 6 io_oeb[23]
port 119 nsew signal output
rlabel metal2 s 97722 199504 97778 200304 6 io_oeb[24]
port 120 nsew signal output
rlabel metal2 s 101678 199504 101734 200304 6 io_oeb[25]
port 121 nsew signal output
rlabel metal2 s 105726 199504 105782 200304 6 io_oeb[26]
port 122 nsew signal output
rlabel metal2 s 109682 199504 109738 200304 6 io_oeb[27]
port 123 nsew signal output
rlabel metal2 s 113638 199504 113694 200304 6 io_oeb[28]
port 124 nsew signal output
rlabel metal2 s 117686 199504 117742 200304 6 io_oeb[29]
port 125 nsew signal output
rlabel metal2 s 9954 199504 10010 200304 6 io_oeb[2]
port 126 nsew signal output
rlabel metal2 s 121642 199504 121698 200304 6 io_oeb[30]
port 127 nsew signal output
rlabel metal2 s 125598 199504 125654 200304 6 io_oeb[31]
port 128 nsew signal output
rlabel metal2 s 129646 199504 129702 200304 6 io_oeb[32]
port 129 nsew signal output
rlabel metal2 s 133602 199504 133658 200304 6 io_oeb[33]
port 130 nsew signal output
rlabel metal2 s 137650 199504 137706 200304 6 io_oeb[34]
port 131 nsew signal output
rlabel metal2 s 141606 199504 141662 200304 6 io_oeb[35]
port 132 nsew signal output
rlabel metal2 s 145562 199504 145618 200304 6 io_oeb[36]
port 133 nsew signal output
rlabel metal2 s 149610 199504 149666 200304 6 io_oeb[37]
port 134 nsew signal output
rlabel metal2 s 13910 199504 13966 200304 6 io_oeb[3]
port 135 nsew signal output
rlabel metal2 s 17866 199504 17922 200304 6 io_oeb[4]
port 136 nsew signal output
rlabel metal2 s 21914 199504 21970 200304 6 io_oeb[5]
port 137 nsew signal output
rlabel metal2 s 25870 199504 25926 200304 6 io_oeb[6]
port 138 nsew signal output
rlabel metal2 s 29918 199504 29974 200304 6 io_oeb[7]
port 139 nsew signal output
rlabel metal2 s 33874 199504 33930 200304 6 io_oeb[8]
port 140 nsew signal output
rlabel metal2 s 37830 199504 37886 200304 6 io_oeb[9]
port 141 nsew signal output
rlabel metal2 s 3238 199504 3294 200304 6 io_out[0]
port 142 nsew signal output
rlabel metal2 s 43166 199504 43222 200304 6 io_out[10]
port 143 nsew signal output
rlabel metal2 s 47122 199504 47178 200304 6 io_out[11]
port 144 nsew signal output
rlabel metal2 s 51170 199504 51226 200304 6 io_out[12]
port 145 nsew signal output
rlabel metal2 s 55126 199504 55182 200304 6 io_out[13]
port 146 nsew signal output
rlabel metal2 s 59174 199504 59230 200304 6 io_out[14]
port 147 nsew signal output
rlabel metal2 s 63130 199504 63186 200304 6 io_out[15]
port 148 nsew signal output
rlabel metal2 s 67086 199504 67142 200304 6 io_out[16]
port 149 nsew signal output
rlabel metal2 s 71134 199504 71190 200304 6 io_out[17]
port 150 nsew signal output
rlabel metal2 s 75090 199504 75146 200304 6 io_out[18]
port 151 nsew signal output
rlabel metal2 s 79046 199504 79102 200304 6 io_out[19]
port 152 nsew signal output
rlabel metal2 s 7286 199504 7342 200304 6 io_out[1]
port 153 nsew signal output
rlabel metal2 s 83094 199504 83150 200304 6 io_out[20]
port 154 nsew signal output
rlabel metal2 s 87050 199504 87106 200304 6 io_out[21]
port 155 nsew signal output
rlabel metal2 s 91098 199504 91154 200304 6 io_out[22]
port 156 nsew signal output
rlabel metal2 s 95054 199504 95110 200304 6 io_out[23]
port 157 nsew signal output
rlabel metal2 s 99010 199504 99066 200304 6 io_out[24]
port 158 nsew signal output
rlabel metal2 s 103058 199504 103114 200304 6 io_out[25]
port 159 nsew signal output
rlabel metal2 s 107014 199504 107070 200304 6 io_out[26]
port 160 nsew signal output
rlabel metal2 s 110970 199504 111026 200304 6 io_out[27]
port 161 nsew signal output
rlabel metal2 s 115018 199504 115074 200304 6 io_out[28]
port 162 nsew signal output
rlabel metal2 s 118974 199504 119030 200304 6 io_out[29]
port 163 nsew signal output
rlabel metal2 s 11242 199504 11298 200304 6 io_out[2]
port 164 nsew signal output
rlabel metal2 s 122930 199504 122986 200304 6 io_out[30]
port 165 nsew signal output
rlabel metal2 s 126978 199504 127034 200304 6 io_out[31]
port 166 nsew signal output
rlabel metal2 s 130934 199504 130990 200304 6 io_out[32]
port 167 nsew signal output
rlabel metal2 s 134982 199504 135038 200304 6 io_out[33]
port 168 nsew signal output
rlabel metal2 s 138938 199504 138994 200304 6 io_out[34]
port 169 nsew signal output
rlabel metal2 s 142894 199504 142950 200304 6 io_out[35]
port 170 nsew signal output
rlabel metal2 s 146942 199504 146998 200304 6 io_out[36]
port 171 nsew signal output
rlabel metal2 s 150898 199504 150954 200304 6 io_out[37]
port 172 nsew signal output
rlabel metal2 s 15290 199504 15346 200304 6 io_out[3]
port 173 nsew signal output
rlabel metal2 s 19246 199504 19302 200304 6 io_out[4]
port 174 nsew signal output
rlabel metal2 s 23202 199504 23258 200304 6 io_out[5]
port 175 nsew signal output
rlabel metal2 s 27250 199504 27306 200304 6 io_out[6]
port 176 nsew signal output
rlabel metal2 s 31206 199504 31262 200304 6 io_out[7]
port 177 nsew signal output
rlabel metal2 s 35162 199504 35218 200304 6 io_out[8]
port 178 nsew signal output
rlabel metal2 s 39210 199504 39266 200304 6 io_out[9]
port 179 nsew signal output
rlabel metal2 s 136086 0 136142 800 6 irq[0]
port 180 nsew signal output
rlabel metal2 s 137282 0 137338 800 6 irq[1]
port 181 nsew signal output
rlabel metal2 s 138570 0 138626 800 6 irq[2]
port 182 nsew signal output
rlabel metal2 s 139858 0 139914 800 6 o_csb0
port 183 nsew signal output
rlabel metal2 s 141146 0 141202 800 6 o_csb0_1
port 184 nsew signal output
rlabel metal3 s 197360 7896 198160 8016 6 o_din0[0]
port 185 nsew signal output
rlabel metal2 s 168010 0 168066 800 6 o_din0[10]
port 186 nsew signal output
rlabel metal3 s 197360 110848 198160 110968 6 o_din0[11]
port 187 nsew signal output
rlabel metal2 s 170586 0 170642 800 6 o_din0[12]
port 188 nsew signal output
rlabel metal3 s 0 116696 800 116816 6 o_din0[13]
port 189 nsew signal output
rlabel metal3 s 197360 121592 198160 121712 6 o_din0[14]
port 190 nsew signal output
rlabel metal2 s 174358 0 174414 800 6 o_din0[15]
port 191 nsew signal output
rlabel metal3 s 0 130976 800 131096 6 o_din0[16]
port 192 nsew signal output
rlabel metal3 s 197360 148656 198160 148776 6 o_din0[17]
port 193 nsew signal output
rlabel metal2 s 175646 0 175702 800 6 o_din0[18]
port 194 nsew signal output
rlabel metal2 s 180154 199504 180210 200304 6 o_din0[19]
port 195 nsew signal output
rlabel metal2 s 145010 0 145066 800 6 o_din0[1]
port 196 nsew signal output
rlabel metal2 s 178222 0 178278 800 6 o_din0[20]
port 197 nsew signal output
rlabel metal3 s 0 169192 800 169312 6 o_din0[21]
port 198 nsew signal output
rlabel metal3 s 197360 154096 198160 154216 6 o_din0[22]
port 199 nsew signal output
rlabel metal3 s 0 173952 800 174072 6 o_din0[23]
port 200 nsew signal output
rlabel metal2 s 184662 0 184718 800 6 o_din0[24]
port 201 nsew signal output
rlabel metal2 s 187146 0 187202 800 6 o_din0[25]
port 202 nsew signal output
rlabel metal3 s 0 183472 800 183592 6 o_din0[26]
port 203 nsew signal output
rlabel metal3 s 0 188232 800 188352 6 o_din0[27]
port 204 nsew signal output
rlabel metal2 s 190826 199504 190882 200304 6 o_din0[28]
port 205 nsew signal output
rlabel metal2 s 194874 0 194930 800 6 o_din0[29]
port 206 nsew signal output
rlabel metal3 s 197360 45840 198160 45960 6 o_din0[2]
port 207 nsew signal output
rlabel metal2 s 196162 0 196218 800 6 o_din0[30]
port 208 nsew signal output
rlabel metal2 s 197450 199504 197506 200304 6 o_din0[31]
port 209 nsew signal output
rlabel metal3 s 197360 67464 198160 67584 6 o_din0[3]
port 210 nsew signal output
rlabel metal2 s 157522 199504 157578 200304 6 o_din0[4]
port 211 nsew signal output
rlabel metal3 s 0 69096 800 69216 6 o_din0[5]
port 212 nsew signal output
rlabel metal3 s 197360 83784 198160 83904 6 o_din0[6]
port 213 nsew signal output
rlabel metal3 s 0 78616 800 78736 6 o_din0[7]
port 214 nsew signal output
rlabel metal3 s 197360 105408 198160 105528 6 o_din0[8]
port 215 nsew signal output
rlabel metal2 s 168194 199504 168250 200304 6 o_din0[9]
port 216 nsew signal output
rlabel metal2 s 153566 199504 153622 200304 6 o_din0_1[0]
port 217 nsew signal output
rlabel metal2 s 166722 0 166778 800 6 o_din0_1[10]
port 218 nsew signal output
rlabel metal3 s 0 97656 800 97776 6 o_din0_1[11]
port 219 nsew signal output
rlabel metal2 s 169298 0 169354 800 6 o_din0_1[12]
port 220 nsew signal output
rlabel metal3 s 0 111936 800 112056 6 o_din0_1[13]
port 221 nsew signal output
rlabel metal2 s 173530 199504 173586 200304 6 o_din0_1[14]
port 222 nsew signal output
rlabel metal2 s 173162 0 173218 800 6 o_din0_1[15]
port 223 nsew signal output
rlabel metal3 s 197360 132472 198160 132592 6 o_din0_1[16]
port 224 nsew signal output
rlabel metal3 s 197360 143352 198160 143472 6 o_din0_1[17]
port 225 nsew signal output
rlabel metal3 s 0 145392 800 145512 6 o_din0_1[18]
port 226 nsew signal output
rlabel metal2 s 176934 0 176990 800 6 o_din0_1[19]
port 227 nsew signal output
rlabel metal2 s 154854 199504 154910 200304 6 o_din0_1[1]
port 228 nsew signal output
rlabel metal3 s 0 164432 800 164552 6 o_din0_1[20]
port 229 nsew signal output
rlabel metal2 s 182822 199504 182878 200304 6 o_din0_1[21]
port 230 nsew signal output
rlabel metal2 s 185490 199504 185546 200304 6 o_din0_1[22]
port 231 nsew signal output
rlabel metal3 s 197360 164976 198160 165096 6 o_din0_1[23]
port 232 nsew signal output
rlabel metal2 s 183374 0 183430 800 6 o_din0_1[24]
port 233 nsew signal output
rlabel metal2 s 185950 0 186006 800 6 o_din0_1[25]
port 234 nsew signal output
rlabel metal2 s 189722 0 189778 800 6 o_din0_1[26]
port 235 nsew signal output
rlabel metal2 s 192298 0 192354 800 6 o_din0_1[27]
port 236 nsew signal output
rlabel metal3 s 197360 186600 198160 186720 6 o_din0_1[28]
port 237 nsew signal output
rlabel metal2 s 192114 199504 192170 200304 6 o_din0_1[29]
port 238 nsew signal output
rlabel metal3 s 197360 40400 198160 40520 6 o_din0_1[2]
port 239 nsew signal output
rlabel metal2 s 194782 199504 194838 200304 6 o_din0_1[30]
port 240 nsew signal output
rlabel metal2 s 196162 199504 196218 200304 6 o_din0_1[31]
port 241 nsew signal output
rlabel metal3 s 0 40400 800 40520 6 o_din0_1[3]
port 242 nsew signal output
rlabel metal2 s 153934 0 153990 800 6 o_din0_1[4]
port 243 nsew signal output
rlabel metal3 s 0 64200 800 64320 6 o_din0_1[5]
port 244 nsew signal output
rlabel metal2 s 160374 0 160430 800 6 o_din0_1[6]
port 245 nsew signal output
rlabel metal3 s 0 73856 800 73976 6 o_din0_1[7]
port 246 nsew signal output
rlabel metal3 s 197360 99968 198160 100088 6 o_din0_1[8]
port 247 nsew signal output
rlabel metal2 s 166906 199504 166962 200304 6 o_din0_1[9]
port 248 nsew signal output
rlabel metal3 s 197360 13336 198160 13456 6 o_waddr0[0]
port 249 nsew signal output
rlabel metal2 s 146298 0 146354 800 6 o_waddr0[1]
port 250 nsew signal output
rlabel metal2 s 148874 0 148930 800 6 o_waddr0[2]
port 251 nsew signal output
rlabel metal2 s 150070 0 150126 800 6 o_waddr0[3]
port 252 nsew signal output
rlabel metal2 s 155222 0 155278 800 6 o_waddr0[4]
port 253 nsew signal output
rlabel metal2 s 156510 0 156566 800 6 o_waddr0[5]
port 254 nsew signal output
rlabel metal2 s 160190 199504 160246 200304 6 o_waddr0[6]
port 255 nsew signal output
rlabel metal2 s 161570 199504 161626 200304 6 o_waddr0[7]
port 256 nsew signal output
rlabel metal2 s 165434 0 165490 800 6 o_waddr0[8]
port 257 nsew signal output
rlabel metal2 s 143722 0 143778 800 6 o_waddr0_1[0]
port 258 nsew signal output
rlabel metal3 s 197360 34960 198160 35080 6 o_waddr0_1[1]
port 259 nsew signal output
rlabel metal3 s 0 30880 800 31000 6 o_waddr0_1[2]
port 260 nsew signal output
rlabel metal3 s 0 45160 800 45280 6 o_waddr0_1[3]
port 261 nsew signal output
rlabel metal3 s 0 54680 800 54800 6 o_waddr0_1[4]
port 262 nsew signal output
rlabel metal3 s 197360 78344 198160 78464 6 o_waddr0_1[5]
port 263 nsew signal output
rlabel metal2 s 161570 0 161626 800 6 o_waddr0_1[6]
port 264 nsew signal output
rlabel metal3 s 197360 94528 198160 94648 6 o_waddr0_1[7]
port 265 nsew signal output
rlabel metal2 s 162858 199504 162914 200304 6 o_waddr0_1[8]
port 266 nsew signal output
rlabel metal3 s 0 7080 800 7200 6 o_web0
port 267 nsew signal output
rlabel metal2 s 142434 0 142490 800 6 o_web0_1
port 268 nsew signal output
rlabel metal3 s 197360 18776 198160 18896 6 o_wmask0[0]
port 269 nsew signal output
rlabel metal3 s 0 21360 800 21480 6 o_wmask0[1]
port 270 nsew signal output
rlabel metal3 s 0 35640 800 35760 6 o_wmask0[2]
port 271 nsew signal output
rlabel metal3 s 197360 72904 198160 73024 6 o_wmask0[3]
port 272 nsew signal output
rlabel metal3 s 197360 24216 198160 24336 6 o_wmask0_1[0]
port 273 nsew signal output
rlabel metal2 s 147586 0 147642 800 6 o_wmask0_1[1]
port 274 nsew signal output
rlabel metal3 s 197360 51280 198160 51400 6 o_wmask0_1[2]
port 275 nsew signal output
rlabel metal2 s 151358 0 151414 800 6 o_wmask0_1[3]
port 276 nsew signal output
rlabel metal3 s 197360 2592 198160 2712 6 rst_i
port 277 nsew signal input
rlabel metal4 s 4208 2128 4528 198064 6 vccd1
port 278 nsew power input
rlabel metal4 s 34928 2128 35248 198064 6 vccd1
port 278 nsew power input
rlabel metal4 s 65648 2128 65968 198064 6 vccd1
port 278 nsew power input
rlabel metal4 s 96368 2128 96688 198064 6 vccd1
port 278 nsew power input
rlabel metal4 s 127088 2128 127408 198064 6 vccd1
port 278 nsew power input
rlabel metal4 s 157808 2128 158128 198064 6 vccd1
port 278 nsew power input
rlabel metal4 s 188528 2128 188848 198064 6 vccd1
port 278 nsew power input
rlabel metal4 s 19568 2128 19888 198064 6 vssd1
port 279 nsew ground input
rlabel metal4 s 50288 2128 50608 198064 6 vssd1
port 279 nsew ground input
rlabel metal4 s 81008 2128 81328 198064 6 vssd1
port 279 nsew ground input
rlabel metal4 s 111728 2128 112048 198064 6 vssd1
port 279 nsew ground input
rlabel metal4 s 142448 2128 142768 198064 6 vssd1
port 279 nsew ground input
rlabel metal4 s 173168 2128 173488 198064 6 vssd1
port 279 nsew ground input
rlabel metal2 s 570 0 626 800 6 wb_clk_i
port 280 nsew signal input
rlabel metal2 s 1766 0 1822 800 6 wb_rst_i
port 281 nsew signal input
rlabel metal2 s 3054 0 3110 800 6 wbs_ack_o
port 282 nsew signal output
rlabel metal2 s 8206 0 8262 800 6 wbs_adr_i[0]
port 283 nsew signal input
rlabel metal2 s 51630 0 51686 800 6 wbs_adr_i[10]
port 284 nsew signal input
rlabel metal2 s 55494 0 55550 800 6 wbs_adr_i[11]
port 285 nsew signal input
rlabel metal2 s 59358 0 59414 800 6 wbs_adr_i[12]
port 286 nsew signal input
rlabel metal2 s 63130 0 63186 800 6 wbs_adr_i[13]
port 287 nsew signal input
rlabel metal2 s 66994 0 67050 800 6 wbs_adr_i[14]
port 288 nsew signal input
rlabel metal2 s 70858 0 70914 800 6 wbs_adr_i[15]
port 289 nsew signal input
rlabel metal2 s 74722 0 74778 800 6 wbs_adr_i[16]
port 290 nsew signal input
rlabel metal2 s 78494 0 78550 800 6 wbs_adr_i[17]
port 291 nsew signal input
rlabel metal2 s 82358 0 82414 800 6 wbs_adr_i[18]
port 292 nsew signal input
rlabel metal2 s 86222 0 86278 800 6 wbs_adr_i[19]
port 293 nsew signal input
rlabel metal2 s 13266 0 13322 800 6 wbs_adr_i[1]
port 294 nsew signal input
rlabel metal2 s 89994 0 90050 800 6 wbs_adr_i[20]
port 295 nsew signal input
rlabel metal2 s 93858 0 93914 800 6 wbs_adr_i[21]
port 296 nsew signal input
rlabel metal2 s 97722 0 97778 800 6 wbs_adr_i[22]
port 297 nsew signal input
rlabel metal2 s 101494 0 101550 800 6 wbs_adr_i[23]
port 298 nsew signal input
rlabel metal2 s 105358 0 105414 800 6 wbs_adr_i[24]
port 299 nsew signal input
rlabel metal2 s 109222 0 109278 800 6 wbs_adr_i[25]
port 300 nsew signal input
rlabel metal2 s 112994 0 113050 800 6 wbs_adr_i[26]
port 301 nsew signal input
rlabel metal2 s 116858 0 116914 800 6 wbs_adr_i[27]
port 302 nsew signal input
rlabel metal2 s 120722 0 120778 800 6 wbs_adr_i[28]
port 303 nsew signal input
rlabel metal2 s 124494 0 124550 800 6 wbs_adr_i[29]
port 304 nsew signal input
rlabel metal2 s 18418 0 18474 800 6 wbs_adr_i[2]
port 305 nsew signal input
rlabel metal2 s 128358 0 128414 800 6 wbs_adr_i[30]
port 306 nsew signal input
rlabel metal2 s 132222 0 132278 800 6 wbs_adr_i[31]
port 307 nsew signal input
rlabel metal2 s 23570 0 23626 800 6 wbs_adr_i[3]
port 308 nsew signal input
rlabel metal2 s 28630 0 28686 800 6 wbs_adr_i[4]
port 309 nsew signal input
rlabel metal2 s 32494 0 32550 800 6 wbs_adr_i[5]
port 310 nsew signal input
rlabel metal2 s 36358 0 36414 800 6 wbs_adr_i[6]
port 311 nsew signal input
rlabel metal2 s 40130 0 40186 800 6 wbs_adr_i[7]
port 312 nsew signal input
rlabel metal2 s 43994 0 44050 800 6 wbs_adr_i[8]
port 313 nsew signal input
rlabel metal2 s 47858 0 47914 800 6 wbs_adr_i[9]
port 314 nsew signal input
rlabel metal2 s 4342 0 4398 800 6 wbs_cyc_i
port 315 nsew signal input
rlabel metal2 s 9494 0 9550 800 6 wbs_dat_i[0]
port 316 nsew signal input
rlabel metal2 s 52918 0 52974 800 6 wbs_dat_i[10]
port 317 nsew signal input
rlabel metal2 s 56782 0 56838 800 6 wbs_dat_i[11]
port 318 nsew signal input
rlabel metal2 s 60646 0 60702 800 6 wbs_dat_i[12]
port 319 nsew signal input
rlabel metal2 s 64418 0 64474 800 6 wbs_dat_i[13]
port 320 nsew signal input
rlabel metal2 s 68282 0 68338 800 6 wbs_dat_i[14]
port 321 nsew signal input
rlabel metal2 s 72146 0 72202 800 6 wbs_dat_i[15]
port 322 nsew signal input
rlabel metal2 s 75918 0 75974 800 6 wbs_dat_i[16]
port 323 nsew signal input
rlabel metal2 s 79782 0 79838 800 6 wbs_dat_i[17]
port 324 nsew signal input
rlabel metal2 s 83646 0 83702 800 6 wbs_dat_i[18]
port 325 nsew signal input
rlabel metal2 s 87418 0 87474 800 6 wbs_dat_i[19]
port 326 nsew signal input
rlabel metal2 s 14554 0 14610 800 6 wbs_dat_i[1]
port 327 nsew signal input
rlabel metal2 s 91282 0 91338 800 6 wbs_dat_i[20]
port 328 nsew signal input
rlabel metal2 s 95146 0 95202 800 6 wbs_dat_i[21]
port 329 nsew signal input
rlabel metal2 s 99010 0 99066 800 6 wbs_dat_i[22]
port 330 nsew signal input
rlabel metal2 s 102782 0 102838 800 6 wbs_dat_i[23]
port 331 nsew signal input
rlabel metal2 s 106646 0 106702 800 6 wbs_dat_i[24]
port 332 nsew signal input
rlabel metal2 s 110510 0 110566 800 6 wbs_dat_i[25]
port 333 nsew signal input
rlabel metal2 s 114282 0 114338 800 6 wbs_dat_i[26]
port 334 nsew signal input
rlabel metal2 s 118146 0 118202 800 6 wbs_dat_i[27]
port 335 nsew signal input
rlabel metal2 s 122010 0 122066 800 6 wbs_dat_i[28]
port 336 nsew signal input
rlabel metal2 s 125782 0 125838 800 6 wbs_dat_i[29]
port 337 nsew signal input
rlabel metal2 s 19706 0 19762 800 6 wbs_dat_i[2]
port 338 nsew signal input
rlabel metal2 s 129646 0 129702 800 6 wbs_dat_i[30]
port 339 nsew signal input
rlabel metal2 s 133510 0 133566 800 6 wbs_dat_i[31]
port 340 nsew signal input
rlabel metal2 s 24858 0 24914 800 6 wbs_dat_i[3]
port 341 nsew signal input
rlabel metal2 s 29918 0 29974 800 6 wbs_dat_i[4]
port 342 nsew signal input
rlabel metal2 s 33782 0 33838 800 6 wbs_dat_i[5]
port 343 nsew signal input
rlabel metal2 s 37646 0 37702 800 6 wbs_dat_i[6]
port 344 nsew signal input
rlabel metal2 s 41418 0 41474 800 6 wbs_dat_i[7]
port 345 nsew signal input
rlabel metal2 s 45282 0 45338 800 6 wbs_dat_i[8]
port 346 nsew signal input
rlabel metal2 s 49146 0 49202 800 6 wbs_dat_i[9]
port 347 nsew signal input
rlabel metal2 s 10782 0 10838 800 6 wbs_dat_o[0]
port 348 nsew signal output
rlabel metal2 s 54206 0 54262 800 6 wbs_dat_o[10]
port 349 nsew signal output
rlabel metal2 s 58070 0 58126 800 6 wbs_dat_o[11]
port 350 nsew signal output
rlabel metal2 s 61934 0 61990 800 6 wbs_dat_o[12]
port 351 nsew signal output
rlabel metal2 s 65706 0 65762 800 6 wbs_dat_o[13]
port 352 nsew signal output
rlabel metal2 s 69570 0 69626 800 6 wbs_dat_o[14]
port 353 nsew signal output
rlabel metal2 s 73434 0 73490 800 6 wbs_dat_o[15]
port 354 nsew signal output
rlabel metal2 s 77206 0 77262 800 6 wbs_dat_o[16]
port 355 nsew signal output
rlabel metal2 s 81070 0 81126 800 6 wbs_dat_o[17]
port 356 nsew signal output
rlabel metal2 s 84934 0 84990 800 6 wbs_dat_o[18]
port 357 nsew signal output
rlabel metal2 s 88706 0 88762 800 6 wbs_dat_o[19]
port 358 nsew signal output
rlabel metal2 s 15842 0 15898 800 6 wbs_dat_o[1]
port 359 nsew signal output
rlabel metal2 s 92570 0 92626 800 6 wbs_dat_o[20]
port 360 nsew signal output
rlabel metal2 s 96434 0 96490 800 6 wbs_dat_o[21]
port 361 nsew signal output
rlabel metal2 s 100206 0 100262 800 6 wbs_dat_o[22]
port 362 nsew signal output
rlabel metal2 s 104070 0 104126 800 6 wbs_dat_o[23]
port 363 nsew signal output
rlabel metal2 s 107934 0 107990 800 6 wbs_dat_o[24]
port 364 nsew signal output
rlabel metal2 s 111798 0 111854 800 6 wbs_dat_o[25]
port 365 nsew signal output
rlabel metal2 s 115570 0 115626 800 6 wbs_dat_o[26]
port 366 nsew signal output
rlabel metal2 s 119434 0 119490 800 6 wbs_dat_o[27]
port 367 nsew signal output
rlabel metal2 s 123298 0 123354 800 6 wbs_dat_o[28]
port 368 nsew signal output
rlabel metal2 s 127070 0 127126 800 6 wbs_dat_o[29]
port 369 nsew signal output
rlabel metal2 s 20994 0 21050 800 6 wbs_dat_o[2]
port 370 nsew signal output
rlabel metal2 s 130934 0 130990 800 6 wbs_dat_o[30]
port 371 nsew signal output
rlabel metal2 s 134798 0 134854 800 6 wbs_dat_o[31]
port 372 nsew signal output
rlabel metal2 s 26054 0 26110 800 6 wbs_dat_o[3]
port 373 nsew signal output
rlabel metal2 s 31206 0 31262 800 6 wbs_dat_o[4]
port 374 nsew signal output
rlabel metal2 s 35070 0 35126 800 6 wbs_dat_o[5]
port 375 nsew signal output
rlabel metal2 s 38842 0 38898 800 6 wbs_dat_o[6]
port 376 nsew signal output
rlabel metal2 s 42706 0 42762 800 6 wbs_dat_o[7]
port 377 nsew signal output
rlabel metal2 s 46570 0 46626 800 6 wbs_dat_o[8]
port 378 nsew signal output
rlabel metal2 s 50342 0 50398 800 6 wbs_dat_o[9]
port 379 nsew signal output
rlabel metal2 s 12070 0 12126 800 6 wbs_sel_i[0]
port 380 nsew signal input
rlabel metal2 s 17130 0 17186 800 6 wbs_sel_i[1]
port 381 nsew signal input
rlabel metal2 s 22282 0 22338 800 6 wbs_sel_i[2]
port 382 nsew signal input
rlabel metal2 s 27342 0 27398 800 6 wbs_sel_i[3]
port 383 nsew signal input
rlabel metal2 s 5630 0 5686 800 6 wbs_stb_i
port 384 nsew signal input
rlabel metal2 s 6918 0 6974 800 6 wbs_we_i
port 385 nsew signal input
<< properties >>
string LEFclass BLOCK
string FIXED_BBOX 0 0 198160 200304
string LEFview TRUE
string GDS_FILE /project/openlane/user_proj/runs/user_proj/results/magic/user_proj.gds
string GDS_END 97319928
string GDS_START 1497704
<< end >>

