magic
tech sky130A
magscale 1 2
timestamp 1645589553
<< obsli1 >>
rect 1104 2159 199151 199121
<< obsm1 >>
rect 1104 484 199350 199436
<< metal2 >>
rect 570 200768 626 201568
rect 1766 200768 1822 201568
rect 3054 200768 3110 201568
rect 4250 200768 4306 201568
rect 5538 200768 5594 201568
rect 6826 200768 6882 201568
rect 8022 200768 8078 201568
rect 9310 200768 9366 201568
rect 10598 200768 10654 201568
rect 11794 200768 11850 201568
rect 13082 200768 13138 201568
rect 14278 200768 14334 201568
rect 15566 200768 15622 201568
rect 16854 200768 16910 201568
rect 18050 200768 18106 201568
rect 19338 200768 19394 201568
rect 20626 200768 20682 201568
rect 21822 200768 21878 201568
rect 23110 200768 23166 201568
rect 24398 200768 24454 201568
rect 25594 200768 25650 201568
rect 26882 200768 26938 201568
rect 28078 200768 28134 201568
rect 29366 200768 29422 201568
rect 30654 200768 30710 201568
rect 31850 200768 31906 201568
rect 33138 200768 33194 201568
rect 34426 200768 34482 201568
rect 35622 200768 35678 201568
rect 36910 200768 36966 201568
rect 38198 200768 38254 201568
rect 39394 200768 39450 201568
rect 40682 200768 40738 201568
rect 41878 200768 41934 201568
rect 43166 200768 43222 201568
rect 44454 200768 44510 201568
rect 45650 200768 45706 201568
rect 46938 200768 46994 201568
rect 48226 200768 48282 201568
rect 49422 200768 49478 201568
rect 50710 200768 50766 201568
rect 51998 200768 52054 201568
rect 53194 200768 53250 201568
rect 54482 200768 54538 201568
rect 55678 200768 55734 201568
rect 56966 200768 57022 201568
rect 58254 200768 58310 201568
rect 59450 200768 59506 201568
rect 60738 200768 60794 201568
rect 62026 200768 62082 201568
rect 63222 200768 63278 201568
rect 64510 200768 64566 201568
rect 65798 200768 65854 201568
rect 66994 200768 67050 201568
rect 68282 200768 68338 201568
rect 69478 200768 69534 201568
rect 70766 200768 70822 201568
rect 72054 200768 72110 201568
rect 73250 200768 73306 201568
rect 74538 200768 74594 201568
rect 75826 200768 75882 201568
rect 77022 200768 77078 201568
rect 78310 200768 78366 201568
rect 79598 200768 79654 201568
rect 80794 200768 80850 201568
rect 82082 200768 82138 201568
rect 83278 200768 83334 201568
rect 84566 200768 84622 201568
rect 85854 200768 85910 201568
rect 87050 200768 87106 201568
rect 88338 200768 88394 201568
rect 89626 200768 89682 201568
rect 90822 200768 90878 201568
rect 92110 200768 92166 201568
rect 93398 200768 93454 201568
rect 94594 200768 94650 201568
rect 95882 200768 95938 201568
rect 97078 200768 97134 201568
rect 98366 200768 98422 201568
rect 99654 200768 99710 201568
rect 100850 200768 100906 201568
rect 102138 200768 102194 201568
rect 103426 200768 103482 201568
rect 104622 200768 104678 201568
rect 105910 200768 105966 201568
rect 107106 200768 107162 201568
rect 108394 200768 108450 201568
rect 109682 200768 109738 201568
rect 110878 200768 110934 201568
rect 112166 200768 112222 201568
rect 113454 200768 113510 201568
rect 114650 200768 114706 201568
rect 115938 200768 115994 201568
rect 117226 200768 117282 201568
rect 118422 200768 118478 201568
rect 119710 200768 119766 201568
rect 120906 200768 120962 201568
rect 122194 200768 122250 201568
rect 123482 200768 123538 201568
rect 124678 200768 124734 201568
rect 125966 200768 126022 201568
rect 127254 200768 127310 201568
rect 128450 200768 128506 201568
rect 129738 200768 129794 201568
rect 131026 200768 131082 201568
rect 132222 200768 132278 201568
rect 133510 200768 133566 201568
rect 134706 200768 134762 201568
rect 135994 200768 136050 201568
rect 137282 200768 137338 201568
rect 138478 200768 138534 201568
rect 139766 200768 139822 201568
rect 141054 200768 141110 201568
rect 142250 200768 142306 201568
rect 143538 200768 143594 201568
rect 144826 200768 144882 201568
rect 146022 200768 146078 201568
rect 147310 200768 147366 201568
rect 148506 200768 148562 201568
rect 149794 200768 149850 201568
rect 151082 200768 151138 201568
rect 152278 200768 152334 201568
rect 153566 200768 153622 201568
rect 154854 200768 154910 201568
rect 156050 200768 156106 201568
rect 157338 200768 157394 201568
rect 158626 200768 158682 201568
rect 159822 200768 159878 201568
rect 161110 200768 161166 201568
rect 162306 200768 162362 201568
rect 163594 200768 163650 201568
rect 164882 200768 164938 201568
rect 166078 200768 166134 201568
rect 167366 200768 167422 201568
rect 168654 200768 168710 201568
rect 169850 200768 169906 201568
rect 171138 200768 171194 201568
rect 172426 200768 172482 201568
rect 173622 200768 173678 201568
rect 174910 200768 174966 201568
rect 176106 200768 176162 201568
rect 177394 200768 177450 201568
rect 178682 200768 178738 201568
rect 179878 200768 179934 201568
rect 181166 200768 181222 201568
rect 182454 200768 182510 201568
rect 183650 200768 183706 201568
rect 184938 200768 184994 201568
rect 186226 200768 186282 201568
rect 187422 200768 187478 201568
rect 188710 200768 188766 201568
rect 189906 200768 189962 201568
rect 191194 200768 191250 201568
rect 192482 200768 192538 201568
rect 193678 200768 193734 201568
rect 194966 200768 195022 201568
rect 196254 200768 196310 201568
rect 197450 200768 197506 201568
rect 198738 200768 198794 201568
rect 662 0 718 800
rect 2042 0 2098 800
rect 3422 0 3478 800
rect 4894 0 4950 800
rect 6274 0 6330 800
rect 7746 0 7802 800
rect 9126 0 9182 800
rect 10598 0 10654 800
rect 11978 0 12034 800
rect 13450 0 13506 800
rect 14830 0 14886 800
rect 16302 0 16358 800
rect 17682 0 17738 800
rect 19154 0 19210 800
rect 20534 0 20590 800
rect 22006 0 22062 800
rect 23386 0 23442 800
rect 24858 0 24914 800
rect 26238 0 26294 800
rect 27710 0 27766 800
rect 29090 0 29146 800
rect 30562 0 30618 800
rect 31942 0 31998 800
rect 33414 0 33470 800
rect 34794 0 34850 800
rect 36266 0 36322 800
rect 37646 0 37702 800
rect 39118 0 39174 800
rect 40498 0 40554 800
rect 41970 0 42026 800
rect 43350 0 43406 800
rect 44822 0 44878 800
rect 46202 0 46258 800
rect 47674 0 47730 800
rect 49054 0 49110 800
rect 50526 0 50582 800
rect 51906 0 51962 800
rect 53286 0 53342 800
rect 54758 0 54814 800
rect 56138 0 56194 800
rect 57610 0 57666 800
rect 58990 0 59046 800
rect 60462 0 60518 800
rect 61842 0 61898 800
rect 63314 0 63370 800
rect 64694 0 64750 800
rect 66166 0 66222 800
rect 67546 0 67602 800
rect 69018 0 69074 800
rect 70398 0 70454 800
rect 71870 0 71926 800
rect 73250 0 73306 800
rect 74722 0 74778 800
rect 76102 0 76158 800
rect 77574 0 77630 800
rect 78954 0 79010 800
rect 80426 0 80482 800
rect 81806 0 81862 800
rect 83278 0 83334 800
rect 84658 0 84714 800
rect 86130 0 86186 800
rect 87510 0 87566 800
rect 88982 0 89038 800
rect 90362 0 90418 800
rect 91834 0 91890 800
rect 93214 0 93270 800
rect 94686 0 94742 800
rect 96066 0 96122 800
rect 97538 0 97594 800
rect 98918 0 98974 800
rect 100390 0 100446 800
rect 101770 0 101826 800
rect 103150 0 103206 800
rect 104622 0 104678 800
rect 106002 0 106058 800
rect 107474 0 107530 800
rect 108854 0 108910 800
rect 110326 0 110382 800
rect 111706 0 111762 800
rect 113178 0 113234 800
rect 114558 0 114614 800
rect 116030 0 116086 800
rect 117410 0 117466 800
rect 118882 0 118938 800
rect 120262 0 120318 800
rect 121734 0 121790 800
rect 123114 0 123170 800
rect 124586 0 124642 800
rect 125966 0 126022 800
rect 127438 0 127494 800
rect 128818 0 128874 800
rect 130290 0 130346 800
rect 131670 0 131726 800
rect 133142 0 133198 800
rect 134522 0 134578 800
rect 135994 0 136050 800
rect 137374 0 137430 800
rect 138846 0 138902 800
rect 140226 0 140282 800
rect 141698 0 141754 800
rect 143078 0 143134 800
rect 144550 0 144606 800
rect 145930 0 145986 800
rect 147402 0 147458 800
rect 148782 0 148838 800
rect 150254 0 150310 800
rect 151634 0 151690 800
rect 153014 0 153070 800
rect 154486 0 154542 800
rect 155866 0 155922 800
rect 157338 0 157394 800
rect 158718 0 158774 800
rect 160190 0 160246 800
rect 161570 0 161626 800
rect 163042 0 163098 800
rect 164422 0 164478 800
rect 165894 0 165950 800
rect 167274 0 167330 800
rect 168746 0 168802 800
rect 170126 0 170182 800
rect 171598 0 171654 800
rect 172978 0 173034 800
rect 174450 0 174506 800
rect 175830 0 175886 800
rect 177302 0 177358 800
rect 178682 0 178738 800
rect 180154 0 180210 800
rect 181534 0 181590 800
rect 183006 0 183062 800
rect 184386 0 184442 800
rect 185858 0 185914 800
rect 187238 0 187294 800
rect 188710 0 188766 800
rect 190090 0 190146 800
rect 191562 0 191618 800
rect 192942 0 192998 800
rect 194414 0 194470 800
rect 195794 0 195850 800
rect 197266 0 197322 800
rect 198646 0 198702 800
<< obsm2 >>
rect 682 200712 1710 200768
rect 1878 200712 2998 200768
rect 3166 200712 4194 200768
rect 4362 200712 5482 200768
rect 5650 200712 6770 200768
rect 6938 200712 7966 200768
rect 8134 200712 9254 200768
rect 9422 200712 10542 200768
rect 10710 200712 11738 200768
rect 11906 200712 13026 200768
rect 13194 200712 14222 200768
rect 14390 200712 15510 200768
rect 15678 200712 16798 200768
rect 16966 200712 17994 200768
rect 18162 200712 19282 200768
rect 19450 200712 20570 200768
rect 20738 200712 21766 200768
rect 21934 200712 23054 200768
rect 23222 200712 24342 200768
rect 24510 200712 25538 200768
rect 25706 200712 26826 200768
rect 26994 200712 28022 200768
rect 28190 200712 29310 200768
rect 29478 200712 30598 200768
rect 30766 200712 31794 200768
rect 31962 200712 33082 200768
rect 33250 200712 34370 200768
rect 34538 200712 35566 200768
rect 35734 200712 36854 200768
rect 37022 200712 38142 200768
rect 38310 200712 39338 200768
rect 39506 200712 40626 200768
rect 40794 200712 41822 200768
rect 41990 200712 43110 200768
rect 43278 200712 44398 200768
rect 44566 200712 45594 200768
rect 45762 200712 46882 200768
rect 47050 200712 48170 200768
rect 48338 200712 49366 200768
rect 49534 200712 50654 200768
rect 50822 200712 51942 200768
rect 52110 200712 53138 200768
rect 53306 200712 54426 200768
rect 54594 200712 55622 200768
rect 55790 200712 56910 200768
rect 57078 200712 58198 200768
rect 58366 200712 59394 200768
rect 59562 200712 60682 200768
rect 60850 200712 61970 200768
rect 62138 200712 63166 200768
rect 63334 200712 64454 200768
rect 64622 200712 65742 200768
rect 65910 200712 66938 200768
rect 67106 200712 68226 200768
rect 68394 200712 69422 200768
rect 69590 200712 70710 200768
rect 70878 200712 71998 200768
rect 72166 200712 73194 200768
rect 73362 200712 74482 200768
rect 74650 200712 75770 200768
rect 75938 200712 76966 200768
rect 77134 200712 78254 200768
rect 78422 200712 79542 200768
rect 79710 200712 80738 200768
rect 80906 200712 82026 200768
rect 82194 200712 83222 200768
rect 83390 200712 84510 200768
rect 84678 200712 85798 200768
rect 85966 200712 86994 200768
rect 87162 200712 88282 200768
rect 88450 200712 89570 200768
rect 89738 200712 90766 200768
rect 90934 200712 92054 200768
rect 92222 200712 93342 200768
rect 93510 200712 94538 200768
rect 94706 200712 95826 200768
rect 95994 200712 97022 200768
rect 97190 200712 98310 200768
rect 98478 200712 99598 200768
rect 99766 200712 100794 200768
rect 100962 200712 102082 200768
rect 102250 200712 103370 200768
rect 103538 200712 104566 200768
rect 104734 200712 105854 200768
rect 106022 200712 107050 200768
rect 107218 200712 108338 200768
rect 108506 200712 109626 200768
rect 109794 200712 110822 200768
rect 110990 200712 112110 200768
rect 112278 200712 113398 200768
rect 113566 200712 114594 200768
rect 114762 200712 115882 200768
rect 116050 200712 117170 200768
rect 117338 200712 118366 200768
rect 118534 200712 119654 200768
rect 119822 200712 120850 200768
rect 121018 200712 122138 200768
rect 122306 200712 123426 200768
rect 123594 200712 124622 200768
rect 124790 200712 125910 200768
rect 126078 200712 127198 200768
rect 127366 200712 128394 200768
rect 128562 200712 129682 200768
rect 129850 200712 130970 200768
rect 131138 200712 132166 200768
rect 132334 200712 133454 200768
rect 133622 200712 134650 200768
rect 134818 200712 135938 200768
rect 136106 200712 137226 200768
rect 137394 200712 138422 200768
rect 138590 200712 139710 200768
rect 139878 200712 140998 200768
rect 141166 200712 142194 200768
rect 142362 200712 143482 200768
rect 143650 200712 144770 200768
rect 144938 200712 145966 200768
rect 146134 200712 147254 200768
rect 147422 200712 148450 200768
rect 148618 200712 149738 200768
rect 149906 200712 151026 200768
rect 151194 200712 152222 200768
rect 152390 200712 153510 200768
rect 153678 200712 154798 200768
rect 154966 200712 155994 200768
rect 156162 200712 157282 200768
rect 157450 200712 158570 200768
rect 158738 200712 159766 200768
rect 159934 200712 161054 200768
rect 161222 200712 162250 200768
rect 162418 200712 163538 200768
rect 163706 200712 164826 200768
rect 164994 200712 166022 200768
rect 166190 200712 167310 200768
rect 167478 200712 168598 200768
rect 168766 200712 169794 200768
rect 169962 200712 171082 200768
rect 171250 200712 172370 200768
rect 172538 200712 173566 200768
rect 173734 200712 174854 200768
rect 175022 200712 176050 200768
rect 176218 200712 177338 200768
rect 177506 200712 178626 200768
rect 178794 200712 179822 200768
rect 179990 200712 181110 200768
rect 181278 200712 182398 200768
rect 182566 200712 183594 200768
rect 183762 200712 184882 200768
rect 185050 200712 186170 200768
rect 186338 200712 187366 200768
rect 187534 200712 188654 200768
rect 188822 200712 189850 200768
rect 190018 200712 191138 200768
rect 191306 200712 192426 200768
rect 192594 200712 193622 200768
rect 193790 200712 194910 200768
rect 195078 200712 196198 200768
rect 196366 200712 197394 200768
rect 197562 200712 198682 200768
rect 198850 200712 199344 200768
rect 676 856 199344 200712
rect 774 31 1986 856
rect 2154 31 3366 856
rect 3534 31 4838 856
rect 5006 31 6218 856
rect 6386 31 7690 856
rect 7858 31 9070 856
rect 9238 31 10542 856
rect 10710 31 11922 856
rect 12090 31 13394 856
rect 13562 31 14774 856
rect 14942 31 16246 856
rect 16414 31 17626 856
rect 17794 31 19098 856
rect 19266 31 20478 856
rect 20646 31 21950 856
rect 22118 31 23330 856
rect 23498 31 24802 856
rect 24970 31 26182 856
rect 26350 31 27654 856
rect 27822 31 29034 856
rect 29202 31 30506 856
rect 30674 31 31886 856
rect 32054 31 33358 856
rect 33526 31 34738 856
rect 34906 31 36210 856
rect 36378 31 37590 856
rect 37758 31 39062 856
rect 39230 31 40442 856
rect 40610 31 41914 856
rect 42082 31 43294 856
rect 43462 31 44766 856
rect 44934 31 46146 856
rect 46314 31 47618 856
rect 47786 31 48998 856
rect 49166 31 50470 856
rect 50638 31 51850 856
rect 52018 31 53230 856
rect 53398 31 54702 856
rect 54870 31 56082 856
rect 56250 31 57554 856
rect 57722 31 58934 856
rect 59102 31 60406 856
rect 60574 31 61786 856
rect 61954 31 63258 856
rect 63426 31 64638 856
rect 64806 31 66110 856
rect 66278 31 67490 856
rect 67658 31 68962 856
rect 69130 31 70342 856
rect 70510 31 71814 856
rect 71982 31 73194 856
rect 73362 31 74666 856
rect 74834 31 76046 856
rect 76214 31 77518 856
rect 77686 31 78898 856
rect 79066 31 80370 856
rect 80538 31 81750 856
rect 81918 31 83222 856
rect 83390 31 84602 856
rect 84770 31 86074 856
rect 86242 31 87454 856
rect 87622 31 88926 856
rect 89094 31 90306 856
rect 90474 31 91778 856
rect 91946 31 93158 856
rect 93326 31 94630 856
rect 94798 31 96010 856
rect 96178 31 97482 856
rect 97650 31 98862 856
rect 99030 31 100334 856
rect 100502 31 101714 856
rect 101882 31 103094 856
rect 103262 31 104566 856
rect 104734 31 105946 856
rect 106114 31 107418 856
rect 107586 31 108798 856
rect 108966 31 110270 856
rect 110438 31 111650 856
rect 111818 31 113122 856
rect 113290 31 114502 856
rect 114670 31 115974 856
rect 116142 31 117354 856
rect 117522 31 118826 856
rect 118994 31 120206 856
rect 120374 31 121678 856
rect 121846 31 123058 856
rect 123226 31 124530 856
rect 124698 31 125910 856
rect 126078 31 127382 856
rect 127550 31 128762 856
rect 128930 31 130234 856
rect 130402 31 131614 856
rect 131782 31 133086 856
rect 133254 31 134466 856
rect 134634 31 135938 856
rect 136106 31 137318 856
rect 137486 31 138790 856
rect 138958 31 140170 856
rect 140338 31 141642 856
rect 141810 31 143022 856
rect 143190 31 144494 856
rect 144662 31 145874 856
rect 146042 31 147346 856
rect 147514 31 148726 856
rect 148894 31 150198 856
rect 150366 31 151578 856
rect 151746 31 152958 856
rect 153126 31 154430 856
rect 154598 31 155810 856
rect 155978 31 157282 856
rect 157450 31 158662 856
rect 158830 31 160134 856
rect 160302 31 161514 856
rect 161682 31 162986 856
rect 163154 31 164366 856
rect 164534 31 165838 856
rect 166006 31 167218 856
rect 167386 31 168690 856
rect 168858 31 170070 856
rect 170238 31 171542 856
rect 171710 31 172922 856
rect 173090 31 174394 856
rect 174562 31 175774 856
rect 175942 31 177246 856
rect 177414 31 178626 856
rect 178794 31 180098 856
rect 180266 31 181478 856
rect 181646 31 182950 856
rect 183118 31 184330 856
rect 184498 31 185802 856
rect 185970 31 187182 856
rect 187350 31 188654 856
rect 188822 31 190034 856
rect 190202 31 191506 856
rect 191674 31 192886 856
rect 193054 31 194358 856
rect 194526 31 195738 856
rect 195906 31 197210 856
rect 197378 31 198590 856
rect 198758 31 199344 856
<< metal3 >>
rect 0 199248 800 199368
rect 198624 198840 199424 198960
rect 0 194896 800 195016
rect 198624 193536 199424 193656
rect 0 190544 800 190664
rect 198624 188232 199424 188352
rect 0 186192 800 186312
rect 198624 182928 199424 183048
rect 0 181704 800 181824
rect 198624 177624 199424 177744
rect 0 177352 800 177472
rect 0 173000 800 173120
rect 198624 172320 199424 172440
rect 0 168648 800 168768
rect 198624 167016 199424 167136
rect 0 164296 800 164416
rect 198624 161712 199424 161832
rect 0 159808 800 159928
rect 198624 156408 199424 156528
rect 0 155456 800 155576
rect 0 151104 800 151224
rect 198624 151104 199424 151224
rect 0 146752 800 146872
rect 198624 145800 199424 145920
rect 0 142264 800 142384
rect 198624 140496 199424 140616
rect 0 137912 800 138032
rect 198624 135192 199424 135312
rect 0 133560 800 133680
rect 198624 129888 199424 130008
rect 0 129208 800 129328
rect 0 124856 800 124976
rect 198624 124584 199424 124704
rect 0 120368 800 120488
rect 198624 119280 199424 119400
rect 0 116016 800 116136
rect 198624 113976 199424 114096
rect 0 111664 800 111784
rect 198624 108672 199424 108792
rect 0 107312 800 107432
rect 198624 103368 199424 103488
rect 0 102960 800 103080
rect 0 98472 800 98592
rect 198624 98064 199424 98184
rect 0 94120 800 94240
rect 198624 92760 199424 92880
rect 0 89768 800 89888
rect 198624 87456 199424 87576
rect 0 85416 800 85536
rect 198624 82152 199424 82272
rect 0 80928 800 81048
rect 198624 76848 199424 76968
rect 0 76576 800 76696
rect 0 72224 800 72344
rect 198624 71544 199424 71664
rect 0 67872 800 67992
rect 198624 66240 199424 66360
rect 0 63520 800 63640
rect 198624 60936 199424 61056
rect 0 59032 800 59152
rect 198624 55632 199424 55752
rect 0 54680 800 54800
rect 0 50328 800 50448
rect 198624 50328 199424 50448
rect 0 45976 800 46096
rect 198624 45024 199424 45144
rect 0 41488 800 41608
rect 198624 39720 199424 39840
rect 0 37136 800 37256
rect 198624 34416 199424 34536
rect 0 32784 800 32904
rect 198624 29112 199424 29232
rect 0 28432 800 28552
rect 0 24080 800 24200
rect 198624 23808 199424 23928
rect 0 19592 800 19712
rect 198624 18504 199424 18624
rect 0 15240 800 15360
rect 198624 13200 199424 13320
rect 0 10888 800 11008
rect 198624 7896 199424 8016
rect 0 6536 800 6656
rect 198624 2592 199424 2712
rect 0 2184 800 2304
<< obsm3 >>
rect 749 199448 199259 199613
rect 880 199168 199259 199448
rect 749 199040 199259 199168
rect 749 198760 198544 199040
rect 749 195096 199259 198760
rect 880 194816 199259 195096
rect 749 193736 199259 194816
rect 749 193456 198544 193736
rect 749 190744 199259 193456
rect 880 190464 199259 190744
rect 749 188432 199259 190464
rect 749 188152 198544 188432
rect 749 186392 199259 188152
rect 880 186112 199259 186392
rect 749 183128 199259 186112
rect 749 182848 198544 183128
rect 749 181904 199259 182848
rect 880 181624 199259 181904
rect 749 177824 199259 181624
rect 749 177552 198544 177824
rect 880 177544 198544 177552
rect 880 177272 199259 177544
rect 749 173200 199259 177272
rect 880 172920 199259 173200
rect 749 172520 199259 172920
rect 749 172240 198544 172520
rect 749 168848 199259 172240
rect 880 168568 199259 168848
rect 749 167216 199259 168568
rect 749 166936 198544 167216
rect 749 164496 199259 166936
rect 880 164216 199259 164496
rect 749 161912 199259 164216
rect 749 161632 198544 161912
rect 749 160008 199259 161632
rect 880 159728 199259 160008
rect 749 156608 199259 159728
rect 749 156328 198544 156608
rect 749 155656 199259 156328
rect 880 155376 199259 155656
rect 749 151304 199259 155376
rect 880 151024 198544 151304
rect 749 146952 199259 151024
rect 880 146672 199259 146952
rect 749 146000 199259 146672
rect 749 145720 198544 146000
rect 749 142464 199259 145720
rect 880 142184 199259 142464
rect 749 140696 199259 142184
rect 749 140416 198544 140696
rect 749 138112 199259 140416
rect 880 137832 199259 138112
rect 749 135392 199259 137832
rect 749 135112 198544 135392
rect 749 133760 199259 135112
rect 880 133480 199259 133760
rect 749 130088 199259 133480
rect 749 129808 198544 130088
rect 749 129408 199259 129808
rect 880 129128 199259 129408
rect 749 125056 199259 129128
rect 880 124784 199259 125056
rect 880 124776 198544 124784
rect 749 124504 198544 124776
rect 749 120568 199259 124504
rect 880 120288 199259 120568
rect 749 119480 199259 120288
rect 749 119200 198544 119480
rect 749 116216 199259 119200
rect 880 115936 199259 116216
rect 749 114176 199259 115936
rect 749 113896 198544 114176
rect 749 111864 199259 113896
rect 880 111584 199259 111864
rect 749 108872 199259 111584
rect 749 108592 198544 108872
rect 749 107512 199259 108592
rect 880 107232 199259 107512
rect 749 103568 199259 107232
rect 749 103288 198544 103568
rect 749 103160 199259 103288
rect 880 102880 199259 103160
rect 749 98672 199259 102880
rect 880 98392 199259 98672
rect 749 98264 199259 98392
rect 749 97984 198544 98264
rect 749 94320 199259 97984
rect 880 94040 199259 94320
rect 749 92960 199259 94040
rect 749 92680 198544 92960
rect 749 89968 199259 92680
rect 880 89688 199259 89968
rect 749 87656 199259 89688
rect 749 87376 198544 87656
rect 749 85616 199259 87376
rect 880 85336 199259 85616
rect 749 82352 199259 85336
rect 749 82072 198544 82352
rect 749 81128 199259 82072
rect 880 80848 199259 81128
rect 749 77048 199259 80848
rect 749 76776 198544 77048
rect 880 76768 198544 76776
rect 880 76496 199259 76768
rect 749 72424 199259 76496
rect 880 72144 199259 72424
rect 749 71744 199259 72144
rect 749 71464 198544 71744
rect 749 68072 199259 71464
rect 880 67792 199259 68072
rect 749 66440 199259 67792
rect 749 66160 198544 66440
rect 749 63720 199259 66160
rect 880 63440 199259 63720
rect 749 61136 199259 63440
rect 749 60856 198544 61136
rect 749 59232 199259 60856
rect 880 58952 199259 59232
rect 749 55832 199259 58952
rect 749 55552 198544 55832
rect 749 54880 199259 55552
rect 880 54600 199259 54880
rect 749 50528 199259 54600
rect 880 50248 198544 50528
rect 749 46176 199259 50248
rect 880 45896 199259 46176
rect 749 45224 199259 45896
rect 749 44944 198544 45224
rect 749 41688 199259 44944
rect 880 41408 199259 41688
rect 749 39920 199259 41408
rect 749 39640 198544 39920
rect 749 37336 199259 39640
rect 880 37056 199259 37336
rect 749 34616 199259 37056
rect 749 34336 198544 34616
rect 749 32984 199259 34336
rect 880 32704 199259 32984
rect 749 29312 199259 32704
rect 749 29032 198544 29312
rect 749 28632 199259 29032
rect 880 28352 199259 28632
rect 749 24280 199259 28352
rect 880 24008 199259 24280
rect 880 24000 198544 24008
rect 749 23728 198544 24000
rect 749 19792 199259 23728
rect 880 19512 199259 19792
rect 749 18704 199259 19512
rect 749 18424 198544 18704
rect 749 15440 199259 18424
rect 880 15160 199259 15440
rect 749 13400 199259 15160
rect 749 13120 198544 13400
rect 749 11088 199259 13120
rect 880 10808 199259 11088
rect 749 8096 199259 10808
rect 749 7816 198544 8096
rect 749 6736 199259 7816
rect 880 6456 199259 6736
rect 749 2792 199259 6456
rect 749 2512 198544 2792
rect 749 2384 199259 2512
rect 880 2104 199259 2384
rect 749 35 199259 2104
<< metal4 >>
rect 4208 2128 4528 199152
rect 19568 2128 19888 199152
rect 34928 2128 35248 199152
rect 50288 2128 50608 199152
rect 65648 2128 65968 199152
rect 81008 2128 81328 199152
rect 96368 2128 96688 199152
rect 111728 2128 112048 199152
rect 127088 2128 127408 199152
rect 142448 2128 142768 199152
rect 157808 2128 158128 199152
rect 173168 2128 173488 199152
rect 188528 2128 188848 199152
<< obsm4 >>
rect 8891 199232 196637 199613
rect 8891 2048 19488 199232
rect 19968 2048 34848 199232
rect 35328 2048 50208 199232
rect 50688 2048 65568 199232
rect 66048 2048 80928 199232
rect 81408 2048 96288 199232
rect 96768 2048 111648 199232
rect 112128 2048 127008 199232
rect 127488 2048 142368 199232
rect 142848 2048 157728 199232
rect 158208 2048 173088 199232
rect 173568 2048 188448 199232
rect 188928 2048 196637 199232
rect 8891 1123 196637 2048
<< labels >>
rlabel metal2 s 155866 0 155922 800 6 clk_i
port 1 nsew signal input
rlabel metal2 s 158718 0 158774 800 6 i_dout0[0]
port 2 nsew signal input
rlabel metal3 s 0 102960 800 103080 6 i_dout0[10]
port 3 nsew signal input
rlabel metal2 s 166078 200768 166134 201568 6 i_dout0[11]
port 4 nsew signal input
rlabel metal2 s 167366 200768 167422 201568 6 i_dout0[12]
port 5 nsew signal input
rlabel metal3 s 0 116016 800 116136 6 i_dout0[13]
port 6 nsew signal input
rlabel metal3 s 198624 98064 199424 98184 6 i_dout0[14]
port 7 nsew signal input
rlabel metal3 s 198624 113976 199424 114096 6 i_dout0[15]
port 8 nsew signal input
rlabel metal3 s 0 124856 800 124976 6 i_dout0[16]
port 9 nsew signal input
rlabel metal3 s 198624 124584 199424 124704 6 i_dout0[17]
port 10 nsew signal input
rlabel metal3 s 0 133560 800 133680 6 i_dout0[18]
port 11 nsew signal input
rlabel metal2 s 178682 200768 178738 201568 6 i_dout0[19]
port 12 nsew signal input
rlabel metal3 s 0 15240 800 15360 6 i_dout0[1]
port 13 nsew signal input
rlabel metal2 s 181166 200768 181222 201568 6 i_dout0[20]
port 14 nsew signal input
rlabel metal2 s 187238 0 187294 800 6 i_dout0[21]
port 15 nsew signal input
rlabel metal3 s 0 159808 800 159928 6 i_dout0[22]
port 16 nsew signal input
rlabel metal2 s 186226 200768 186282 201568 6 i_dout0[23]
port 17 nsew signal input
rlabel metal3 s 198624 172320 199424 172440 6 i_dout0[24]
port 18 nsew signal input
rlabel metal2 s 188710 200768 188766 201568 6 i_dout0[25]
port 19 nsew signal input
rlabel metal3 s 0 173000 800 173120 6 i_dout0[26]
port 20 nsew signal input
rlabel metal3 s 0 177352 800 177472 6 i_dout0[27]
port 21 nsew signal input
rlabel metal3 s 198624 188232 199424 188352 6 i_dout0[28]
port 22 nsew signal input
rlabel metal2 s 198646 0 198702 800 6 i_dout0[29]
port 23 nsew signal input
rlabel metal3 s 198624 34416 199424 34536 6 i_dout0[2]
port 24 nsew signal input
rlabel metal3 s 0 194896 800 195016 6 i_dout0[30]
port 25 nsew signal input
rlabel metal3 s 198624 198840 199424 198960 6 i_dout0[31]
port 26 nsew signal input
rlabel metal3 s 198624 50328 199424 50448 6 i_dout0[3]
port 27 nsew signal input
rlabel metal3 s 198624 66240 199424 66360 6 i_dout0[4]
port 28 nsew signal input
rlabel metal2 s 154854 200768 154910 201568 6 i_dout0[5]
port 29 nsew signal input
rlabel metal3 s 0 72224 800 72344 6 i_dout0[6]
port 30 nsew signal input
rlabel metal2 s 170126 0 170182 800 6 i_dout0[7]
port 31 nsew signal input
rlabel metal2 s 161110 200768 161166 201568 6 i_dout0[8]
port 32 nsew signal input
rlabel metal2 s 178682 0 178738 800 6 i_dout0[9]
port 33 nsew signal input
rlabel metal2 s 160190 0 160246 800 6 i_dout0_1[0]
port 34 nsew signal input
rlabel metal3 s 198624 87456 199424 87576 6 i_dout0_1[10]
port 35 nsew signal input
rlabel metal3 s 0 107312 800 107432 6 i_dout0_1[11]
port 36 nsew signal input
rlabel metal2 s 183006 0 183062 800 6 i_dout0_1[12]
port 37 nsew signal input
rlabel metal2 s 168654 200768 168710 201568 6 i_dout0_1[13]
port 38 nsew signal input
rlabel metal2 s 185858 0 185914 800 6 i_dout0_1[14]
port 39 nsew signal input
rlabel metal3 s 198624 108672 199424 108792 6 i_dout0_1[15]
port 40 nsew signal input
rlabel metal3 s 0 120368 800 120488 6 i_dout0_1[16]
port 41 nsew signal input
rlabel metal3 s 0 129208 800 129328 6 i_dout0_1[17]
port 42 nsew signal input
rlabel metal2 s 177394 200768 177450 201568 6 i_dout0_1[18]
port 43 nsew signal input
rlabel metal3 s 198624 135192 199424 135312 6 i_dout0_1[19]
port 44 nsew signal input
rlabel metal2 s 161570 0 161626 800 6 i_dout0_1[1]
port 45 nsew signal input
rlabel metal3 s 198624 140496 199424 140616 6 i_dout0_1[20]
port 46 nsew signal input
rlabel metal3 s 0 155456 800 155576 6 i_dout0_1[21]
port 47 nsew signal input
rlabel metal2 s 183650 200768 183706 201568 6 i_dout0_1[22]
port 48 nsew signal input
rlabel metal3 s 198624 156408 199424 156528 6 i_dout0_1[23]
port 49 nsew signal input
rlabel metal3 s 198624 167016 199424 167136 6 i_dout0_1[24]
port 50 nsew signal input
rlabel metal2 s 190090 0 190146 800 6 i_dout0_1[25]
port 51 nsew signal input
rlabel metal2 s 191562 0 191618 800 6 i_dout0_1[26]
port 52 nsew signal input
rlabel metal3 s 198624 182928 199424 183048 6 i_dout0_1[27]
port 53 nsew signal input
rlabel metal2 s 195794 0 195850 800 6 i_dout0_1[28]
port 54 nsew signal input
rlabel metal3 s 0 186192 800 186312 6 i_dout0_1[29]
port 55 nsew signal input
rlabel metal2 s 163042 0 163098 800 6 i_dout0_1[2]
port 56 nsew signal input
rlabel metal3 s 0 190544 800 190664 6 i_dout0_1[30]
port 57 nsew signal input
rlabel metal2 s 197450 200768 197506 201568 6 i_dout0_1[31]
port 58 nsew signal input
rlabel metal2 s 165894 0 165950 800 6 i_dout0_1[3]
port 59 nsew signal input
rlabel metal2 s 151082 200768 151138 201568 6 i_dout0_1[4]
port 60 nsew signal input
rlabel metal3 s 0 54680 800 54800 6 i_dout0_1[5]
port 61 nsew signal input
rlabel metal3 s 0 67872 800 67992 6 i_dout0_1[6]
port 62 nsew signal input
rlabel metal2 s 159822 200768 159878 201568 6 i_dout0_1[7]
port 63 nsew signal input
rlabel metal3 s 0 89768 800 89888 6 i_dout0_1[8]
port 64 nsew signal input
rlabel metal2 s 177302 0 177358 800 6 i_dout0_1[9]
port 65 nsew signal input
rlabel metal2 s 570 200768 626 201568 6 io_in[0]
port 66 nsew signal input
rlabel metal2 s 38198 200768 38254 201568 6 io_in[10]
port 67 nsew signal input
rlabel metal2 s 41878 200768 41934 201568 6 io_in[11]
port 68 nsew signal input
rlabel metal2 s 45650 200768 45706 201568 6 io_in[12]
port 69 nsew signal input
rlabel metal2 s 49422 200768 49478 201568 6 io_in[13]
port 70 nsew signal input
rlabel metal2 s 53194 200768 53250 201568 6 io_in[14]
port 71 nsew signal input
rlabel metal2 s 56966 200768 57022 201568 6 io_in[15]
port 72 nsew signal input
rlabel metal2 s 60738 200768 60794 201568 6 io_in[16]
port 73 nsew signal input
rlabel metal2 s 64510 200768 64566 201568 6 io_in[17]
port 74 nsew signal input
rlabel metal2 s 68282 200768 68338 201568 6 io_in[18]
port 75 nsew signal input
rlabel metal2 s 72054 200768 72110 201568 6 io_in[19]
port 76 nsew signal input
rlabel metal2 s 4250 200768 4306 201568 6 io_in[1]
port 77 nsew signal input
rlabel metal2 s 75826 200768 75882 201568 6 io_in[20]
port 78 nsew signal input
rlabel metal2 s 79598 200768 79654 201568 6 io_in[21]
port 79 nsew signal input
rlabel metal2 s 83278 200768 83334 201568 6 io_in[22]
port 80 nsew signal input
rlabel metal2 s 87050 200768 87106 201568 6 io_in[23]
port 81 nsew signal input
rlabel metal2 s 90822 200768 90878 201568 6 io_in[24]
port 82 nsew signal input
rlabel metal2 s 94594 200768 94650 201568 6 io_in[25]
port 83 nsew signal input
rlabel metal2 s 98366 200768 98422 201568 6 io_in[26]
port 84 nsew signal input
rlabel metal2 s 102138 200768 102194 201568 6 io_in[27]
port 85 nsew signal input
rlabel metal2 s 105910 200768 105966 201568 6 io_in[28]
port 86 nsew signal input
rlabel metal2 s 109682 200768 109738 201568 6 io_in[29]
port 87 nsew signal input
rlabel metal2 s 8022 200768 8078 201568 6 io_in[2]
port 88 nsew signal input
rlabel metal2 s 113454 200768 113510 201568 6 io_in[30]
port 89 nsew signal input
rlabel metal2 s 117226 200768 117282 201568 6 io_in[31]
port 90 nsew signal input
rlabel metal2 s 120906 200768 120962 201568 6 io_in[32]
port 91 nsew signal input
rlabel metal2 s 124678 200768 124734 201568 6 io_in[33]
port 92 nsew signal input
rlabel metal2 s 128450 200768 128506 201568 6 io_in[34]
port 93 nsew signal input
rlabel metal2 s 132222 200768 132278 201568 6 io_in[35]
port 94 nsew signal input
rlabel metal2 s 135994 200768 136050 201568 6 io_in[36]
port 95 nsew signal input
rlabel metal2 s 139766 200768 139822 201568 6 io_in[37]
port 96 nsew signal input
rlabel metal2 s 11794 200768 11850 201568 6 io_in[3]
port 97 nsew signal input
rlabel metal2 s 15566 200768 15622 201568 6 io_in[4]
port 98 nsew signal input
rlabel metal2 s 19338 200768 19394 201568 6 io_in[5]
port 99 nsew signal input
rlabel metal2 s 23110 200768 23166 201568 6 io_in[6]
port 100 nsew signal input
rlabel metal2 s 26882 200768 26938 201568 6 io_in[7]
port 101 nsew signal input
rlabel metal2 s 30654 200768 30710 201568 6 io_in[8]
port 102 nsew signal input
rlabel metal2 s 34426 200768 34482 201568 6 io_in[9]
port 103 nsew signal input
rlabel metal2 s 1766 200768 1822 201568 6 io_oeb[0]
port 104 nsew signal output
rlabel metal2 s 39394 200768 39450 201568 6 io_oeb[10]
port 105 nsew signal output
rlabel metal2 s 43166 200768 43222 201568 6 io_oeb[11]
port 106 nsew signal output
rlabel metal2 s 46938 200768 46994 201568 6 io_oeb[12]
port 107 nsew signal output
rlabel metal2 s 50710 200768 50766 201568 6 io_oeb[13]
port 108 nsew signal output
rlabel metal2 s 54482 200768 54538 201568 6 io_oeb[14]
port 109 nsew signal output
rlabel metal2 s 58254 200768 58310 201568 6 io_oeb[15]
port 110 nsew signal output
rlabel metal2 s 62026 200768 62082 201568 6 io_oeb[16]
port 111 nsew signal output
rlabel metal2 s 65798 200768 65854 201568 6 io_oeb[17]
port 112 nsew signal output
rlabel metal2 s 69478 200768 69534 201568 6 io_oeb[18]
port 113 nsew signal output
rlabel metal2 s 73250 200768 73306 201568 6 io_oeb[19]
port 114 nsew signal output
rlabel metal2 s 5538 200768 5594 201568 6 io_oeb[1]
port 115 nsew signal output
rlabel metal2 s 77022 200768 77078 201568 6 io_oeb[20]
port 116 nsew signal output
rlabel metal2 s 80794 200768 80850 201568 6 io_oeb[21]
port 117 nsew signal output
rlabel metal2 s 84566 200768 84622 201568 6 io_oeb[22]
port 118 nsew signal output
rlabel metal2 s 88338 200768 88394 201568 6 io_oeb[23]
port 119 nsew signal output
rlabel metal2 s 92110 200768 92166 201568 6 io_oeb[24]
port 120 nsew signal output
rlabel metal2 s 95882 200768 95938 201568 6 io_oeb[25]
port 121 nsew signal output
rlabel metal2 s 99654 200768 99710 201568 6 io_oeb[26]
port 122 nsew signal output
rlabel metal2 s 103426 200768 103482 201568 6 io_oeb[27]
port 123 nsew signal output
rlabel metal2 s 107106 200768 107162 201568 6 io_oeb[28]
port 124 nsew signal output
rlabel metal2 s 110878 200768 110934 201568 6 io_oeb[29]
port 125 nsew signal output
rlabel metal2 s 9310 200768 9366 201568 6 io_oeb[2]
port 126 nsew signal output
rlabel metal2 s 114650 200768 114706 201568 6 io_oeb[30]
port 127 nsew signal output
rlabel metal2 s 118422 200768 118478 201568 6 io_oeb[31]
port 128 nsew signal output
rlabel metal2 s 122194 200768 122250 201568 6 io_oeb[32]
port 129 nsew signal output
rlabel metal2 s 125966 200768 126022 201568 6 io_oeb[33]
port 130 nsew signal output
rlabel metal2 s 129738 200768 129794 201568 6 io_oeb[34]
port 131 nsew signal output
rlabel metal2 s 133510 200768 133566 201568 6 io_oeb[35]
port 132 nsew signal output
rlabel metal2 s 137282 200768 137338 201568 6 io_oeb[36]
port 133 nsew signal output
rlabel metal2 s 141054 200768 141110 201568 6 io_oeb[37]
port 134 nsew signal output
rlabel metal2 s 13082 200768 13138 201568 6 io_oeb[3]
port 135 nsew signal output
rlabel metal2 s 16854 200768 16910 201568 6 io_oeb[4]
port 136 nsew signal output
rlabel metal2 s 20626 200768 20682 201568 6 io_oeb[5]
port 137 nsew signal output
rlabel metal2 s 24398 200768 24454 201568 6 io_oeb[6]
port 138 nsew signal output
rlabel metal2 s 28078 200768 28134 201568 6 io_oeb[7]
port 139 nsew signal output
rlabel metal2 s 31850 200768 31906 201568 6 io_oeb[8]
port 140 nsew signal output
rlabel metal2 s 35622 200768 35678 201568 6 io_oeb[9]
port 141 nsew signal output
rlabel metal2 s 3054 200768 3110 201568 6 io_out[0]
port 142 nsew signal output
rlabel metal2 s 40682 200768 40738 201568 6 io_out[10]
port 143 nsew signal output
rlabel metal2 s 44454 200768 44510 201568 6 io_out[11]
port 144 nsew signal output
rlabel metal2 s 48226 200768 48282 201568 6 io_out[12]
port 145 nsew signal output
rlabel metal2 s 51998 200768 52054 201568 6 io_out[13]
port 146 nsew signal output
rlabel metal2 s 55678 200768 55734 201568 6 io_out[14]
port 147 nsew signal output
rlabel metal2 s 59450 200768 59506 201568 6 io_out[15]
port 148 nsew signal output
rlabel metal2 s 63222 200768 63278 201568 6 io_out[16]
port 149 nsew signal output
rlabel metal2 s 66994 200768 67050 201568 6 io_out[17]
port 150 nsew signal output
rlabel metal2 s 70766 200768 70822 201568 6 io_out[18]
port 151 nsew signal output
rlabel metal2 s 74538 200768 74594 201568 6 io_out[19]
port 152 nsew signal output
rlabel metal2 s 6826 200768 6882 201568 6 io_out[1]
port 153 nsew signal output
rlabel metal2 s 78310 200768 78366 201568 6 io_out[20]
port 154 nsew signal output
rlabel metal2 s 82082 200768 82138 201568 6 io_out[21]
port 155 nsew signal output
rlabel metal2 s 85854 200768 85910 201568 6 io_out[22]
port 156 nsew signal output
rlabel metal2 s 89626 200768 89682 201568 6 io_out[23]
port 157 nsew signal output
rlabel metal2 s 93398 200768 93454 201568 6 io_out[24]
port 158 nsew signal output
rlabel metal2 s 97078 200768 97134 201568 6 io_out[25]
port 159 nsew signal output
rlabel metal2 s 100850 200768 100906 201568 6 io_out[26]
port 160 nsew signal output
rlabel metal2 s 104622 200768 104678 201568 6 io_out[27]
port 161 nsew signal output
rlabel metal2 s 108394 200768 108450 201568 6 io_out[28]
port 162 nsew signal output
rlabel metal2 s 112166 200768 112222 201568 6 io_out[29]
port 163 nsew signal output
rlabel metal2 s 10598 200768 10654 201568 6 io_out[2]
port 164 nsew signal output
rlabel metal2 s 115938 200768 115994 201568 6 io_out[30]
port 165 nsew signal output
rlabel metal2 s 119710 200768 119766 201568 6 io_out[31]
port 166 nsew signal output
rlabel metal2 s 123482 200768 123538 201568 6 io_out[32]
port 167 nsew signal output
rlabel metal2 s 127254 200768 127310 201568 6 io_out[33]
port 168 nsew signal output
rlabel metal2 s 131026 200768 131082 201568 6 io_out[34]
port 169 nsew signal output
rlabel metal2 s 134706 200768 134762 201568 6 io_out[35]
port 170 nsew signal output
rlabel metal2 s 138478 200768 138534 201568 6 io_out[36]
port 171 nsew signal output
rlabel metal2 s 142250 200768 142306 201568 6 io_out[37]
port 172 nsew signal output
rlabel metal2 s 14278 200768 14334 201568 6 io_out[3]
port 173 nsew signal output
rlabel metal2 s 18050 200768 18106 201568 6 io_out[4]
port 174 nsew signal output
rlabel metal2 s 21822 200768 21878 201568 6 io_out[5]
port 175 nsew signal output
rlabel metal2 s 25594 200768 25650 201568 6 io_out[6]
port 176 nsew signal output
rlabel metal2 s 29366 200768 29422 201568 6 io_out[7]
port 177 nsew signal output
rlabel metal2 s 33138 200768 33194 201568 6 io_out[8]
port 178 nsew signal output
rlabel metal2 s 36910 200768 36966 201568 6 io_out[9]
port 179 nsew signal output
rlabel metal2 s 151634 0 151690 800 6 irq[0]
port 180 nsew signal output
rlabel metal2 s 153014 0 153070 800 6 irq[1]
port 181 nsew signal output
rlabel metal2 s 154486 0 154542 800 6 irq[2]
port 182 nsew signal output
rlabel metal3 s 0 2184 800 2304 6 o_csb0
port 183 nsew signal output
rlabel metal3 s 0 6536 800 6656 6 o_csb0_1
port 184 nsew signal output
rlabel metal3 s 198624 2592 199424 2712 6 o_din0[0]
port 185 nsew signal output
rlabel metal2 s 164882 200768 164938 201568 6 o_din0[10]
port 186 nsew signal output
rlabel metal2 s 181534 0 181590 800 6 o_din0[11]
port 187 nsew signal output
rlabel metal3 s 198624 92760 199424 92880 6 o_din0[12]
port 188 nsew signal output
rlabel metal2 s 184386 0 184442 800 6 o_din0[13]
port 189 nsew signal output
rlabel metal3 s 198624 103368 199424 103488 6 o_din0[14]
port 190 nsew signal output
rlabel metal2 s 173622 200768 173678 201568 6 o_din0[15]
port 191 nsew signal output
rlabel metal3 s 198624 119280 199424 119400 6 o_din0[16]
port 192 nsew signal output
rlabel metal3 s 198624 129888 199424 130008 6 o_din0[17]
port 193 nsew signal output
rlabel metal3 s 0 142264 800 142384 6 o_din0[18]
port 194 nsew signal output
rlabel metal2 s 179878 200768 179934 201568 6 o_din0[19]
port 195 nsew signal output
rlabel metal3 s 198624 18504 199424 18624 6 o_din0[1]
port 196 nsew signal output
rlabel metal2 s 182454 200768 182510 201568 6 o_din0[20]
port 197 nsew signal output
rlabel metal3 s 198624 151104 199424 151224 6 o_din0[21]
port 198 nsew signal output
rlabel metal3 s 0 164296 800 164416 6 o_din0[22]
port 199 nsew signal output
rlabel metal2 s 187422 200768 187478 201568 6 o_din0[23]
port 200 nsew signal output
rlabel metal2 s 188710 0 188766 800 6 o_din0[24]
port 201 nsew signal output
rlabel metal3 s 0 168648 800 168768 6 o_din0[25]
port 202 nsew signal output
rlabel metal2 s 191194 200768 191250 201568 6 o_din0[26]
port 203 nsew signal output
rlabel metal2 s 192482 200768 192538 201568 6 o_din0[27]
port 204 nsew signal output
rlabel metal2 s 197266 0 197322 800 6 o_din0[28]
port 205 nsew signal output
rlabel metal2 s 194966 200768 195022 201568 6 o_din0[29]
port 206 nsew signal output
rlabel metal3 s 0 32784 800 32904 6 o_din0[2]
port 207 nsew signal output
rlabel metal2 s 196254 200768 196310 201568 6 o_din0[30]
port 208 nsew signal output
rlabel metal3 s 0 199248 800 199368 6 o_din0[31]
port 209 nsew signal output
rlabel metal3 s 0 41488 800 41608 6 o_din0[3]
port 210 nsew signal output
rlabel metal3 s 198624 71544 199424 71664 6 o_din0[4]
port 211 nsew signal output
rlabel metal3 s 0 63520 800 63640 6 o_din0[5]
port 212 nsew signal output
rlabel metal3 s 0 80928 800 81048 6 o_din0[6]
port 213 nsew signal output
rlabel metal3 s 0 85416 800 85536 6 o_din0[7]
port 214 nsew signal output
rlabel metal2 s 174450 0 174506 800 6 o_din0[8]
port 215 nsew signal output
rlabel metal3 s 198624 82152 199424 82272 6 o_din0[9]
port 216 nsew signal output
rlabel metal2 s 146022 200768 146078 201568 6 o_din0_1[0]
port 217 nsew signal output
rlabel metal2 s 163594 200768 163650 201568 6 o_din0_1[10]
port 218 nsew signal output
rlabel metal2 s 180154 0 180210 800 6 o_din0_1[11]
port 219 nsew signal output
rlabel metal3 s 0 111664 800 111784 6 o_din0_1[12]
port 220 nsew signal output
rlabel metal2 s 169850 200768 169906 201568 6 o_din0_1[13]
port 221 nsew signal output
rlabel metal2 s 171138 200768 171194 201568 6 o_din0_1[14]
port 222 nsew signal output
rlabel metal2 s 172426 200768 172482 201568 6 o_din0_1[15]
port 223 nsew signal output
rlabel metal2 s 174910 200768 174966 201568 6 o_din0_1[16]
port 224 nsew signal output
rlabel metal2 s 176106 200768 176162 201568 6 o_din0_1[17]
port 225 nsew signal output
rlabel metal3 s 0 137912 800 138032 6 o_din0_1[18]
port 226 nsew signal output
rlabel metal3 s 0 146752 800 146872 6 o_din0_1[19]
port 227 nsew signal output
rlabel metal2 s 148506 200768 148562 201568 6 o_din0_1[1]
port 228 nsew signal output
rlabel metal3 s 0 151104 800 151224 6 o_din0_1[20]
port 229 nsew signal output
rlabel metal3 s 198624 145800 199424 145920 6 o_din0_1[21]
port 230 nsew signal output
rlabel metal2 s 184938 200768 184994 201568 6 o_din0_1[22]
port 231 nsew signal output
rlabel metal3 s 198624 161712 199424 161832 6 o_din0_1[23]
port 232 nsew signal output
rlabel metal3 s 198624 177624 199424 177744 6 o_din0_1[24]
port 233 nsew signal output
rlabel metal2 s 189906 200768 189962 201568 6 o_din0_1[25]
port 234 nsew signal output
rlabel metal2 s 192942 0 192998 800 6 o_din0_1[26]
port 235 nsew signal output
rlabel metal2 s 194414 0 194470 800 6 o_din0_1[27]
port 236 nsew signal output
rlabel metal3 s 0 181704 800 181824 6 o_din0_1[28]
port 237 nsew signal output
rlabel metal2 s 193678 200768 193734 201568 6 o_din0_1[29]
port 238 nsew signal output
rlabel metal3 s 0 28432 800 28552 6 o_din0_1[2]
port 239 nsew signal output
rlabel metal3 s 198624 193536 199424 193656 6 o_din0_1[30]
port 240 nsew signal output
rlabel metal2 s 198738 200768 198794 201568 6 o_din0_1[31]
port 241 nsew signal output
rlabel metal2 s 167274 0 167330 800 6 o_din0_1[3]
port 242 nsew signal output
rlabel metal3 s 0 50328 800 50448 6 o_din0_1[4]
port 243 nsew signal output
rlabel metal3 s 0 59032 800 59152 6 o_din0_1[5]
port 244 nsew signal output
rlabel metal3 s 0 76576 800 76696 6 o_din0_1[6]
port 245 nsew signal output
rlabel metal2 s 171598 0 171654 800 6 o_din0_1[7]
port 246 nsew signal output
rlabel metal2 s 162306 200768 162362 201568 6 o_din0_1[8]
port 247 nsew signal output
rlabel metal3 s 0 98472 800 98592 6 o_din0_1[9]
port 248 nsew signal output
rlabel metal3 s 198624 7896 199424 8016 6 o_waddr0[0]
port 249 nsew signal output
rlabel metal3 s 198624 29112 199424 29232 6 o_waddr0[1]
port 250 nsew signal output
rlabel metal3 s 198624 45024 199424 45144 6 o_waddr0[2]
port 251 nsew signal output
rlabel metal2 s 149794 200768 149850 201568 6 o_waddr0[3]
port 252 nsew signal output
rlabel metal2 s 153566 200768 153622 201568 6 o_waddr0[4]
port 253 nsew signal output
rlabel metal2 s 156050 200768 156106 201568 6 o_waddr0[5]
port 254 nsew signal output
rlabel metal2 s 158626 200768 158682 201568 6 o_waddr0[6]
port 255 nsew signal output
rlabel metal2 s 172978 0 173034 800 6 o_waddr0[7]
port 256 nsew signal output
rlabel metal2 s 175830 0 175886 800 6 o_waddr0[8]
port 257 nsew signal output
rlabel metal3 s 0 10888 800 11008 6 o_waddr0_1[0]
port 258 nsew signal output
rlabel metal3 s 198624 23808 199424 23928 6 o_waddr0_1[1]
port 259 nsew signal output
rlabel metal3 s 198624 39720 199424 39840 6 o_waddr0_1[2]
port 260 nsew signal output
rlabel metal3 s 198624 55632 199424 55752 6 o_waddr0_1[3]
port 261 nsew signal output
rlabel metal2 s 152278 200768 152334 201568 6 o_waddr0_1[4]
port 262 nsew signal output
rlabel metal2 s 168746 0 168802 800 6 o_waddr0_1[5]
port 263 nsew signal output
rlabel metal2 s 157338 200768 157394 201568 6 o_waddr0_1[6]
port 264 nsew signal output
rlabel metal3 s 198624 76848 199424 76968 6 o_waddr0_1[7]
port 265 nsew signal output
rlabel metal3 s 0 94120 800 94240 6 o_waddr0_1[8]
port 266 nsew signal output
rlabel metal2 s 157338 0 157394 800 6 o_web0
port 267 nsew signal output
rlabel metal2 s 143538 200768 143594 201568 6 o_web0_1
port 268 nsew signal output
rlabel metal2 s 147310 200768 147366 201568 6 o_wmask0[0]
port 269 nsew signal output
rlabel metal3 s 0 24080 800 24200 6 o_wmask0[1]
port 270 nsew signal output
rlabel metal2 s 164422 0 164478 800 6 o_wmask0[2]
port 271 nsew signal output
rlabel metal3 s 198624 60936 199424 61056 6 o_wmask0[3]
port 272 nsew signal output
rlabel metal3 s 198624 13200 199424 13320 6 o_wmask0_1[0]
port 273 nsew signal output
rlabel metal3 s 0 19592 800 19712 6 o_wmask0_1[1]
port 274 nsew signal output
rlabel metal3 s 0 37136 800 37256 6 o_wmask0_1[2]
port 275 nsew signal output
rlabel metal3 s 0 45976 800 46096 6 o_wmask0_1[3]
port 276 nsew signal output
rlabel metal2 s 144826 200768 144882 201568 6 rst_i
port 277 nsew signal input
rlabel metal4 s 4208 2128 4528 199152 6 vccd1
port 278 nsew power input
rlabel metal4 s 34928 2128 35248 199152 6 vccd1
port 278 nsew power input
rlabel metal4 s 65648 2128 65968 199152 6 vccd1
port 278 nsew power input
rlabel metal4 s 96368 2128 96688 199152 6 vccd1
port 278 nsew power input
rlabel metal4 s 127088 2128 127408 199152 6 vccd1
port 278 nsew power input
rlabel metal4 s 157808 2128 158128 199152 6 vccd1
port 278 nsew power input
rlabel metal4 s 188528 2128 188848 199152 6 vccd1
port 278 nsew power input
rlabel metal4 s 19568 2128 19888 199152 6 vssd1
port 279 nsew ground input
rlabel metal4 s 50288 2128 50608 199152 6 vssd1
port 279 nsew ground input
rlabel metal4 s 81008 2128 81328 199152 6 vssd1
port 279 nsew ground input
rlabel metal4 s 111728 2128 112048 199152 6 vssd1
port 279 nsew ground input
rlabel metal4 s 142448 2128 142768 199152 6 vssd1
port 279 nsew ground input
rlabel metal4 s 173168 2128 173488 199152 6 vssd1
port 279 nsew ground input
rlabel metal2 s 662 0 718 800 6 wb_clk_i
port 280 nsew signal input
rlabel metal2 s 2042 0 2098 800 6 wb_rst_i
port 281 nsew signal input
rlabel metal2 s 3422 0 3478 800 6 wbs_ack_o
port 282 nsew signal output
rlabel metal2 s 9126 0 9182 800 6 wbs_adr_i[0]
port 283 nsew signal input
rlabel metal2 s 57610 0 57666 800 6 wbs_adr_i[10]
port 284 nsew signal input
rlabel metal2 s 61842 0 61898 800 6 wbs_adr_i[11]
port 285 nsew signal input
rlabel metal2 s 66166 0 66222 800 6 wbs_adr_i[12]
port 286 nsew signal input
rlabel metal2 s 70398 0 70454 800 6 wbs_adr_i[13]
port 287 nsew signal input
rlabel metal2 s 74722 0 74778 800 6 wbs_adr_i[14]
port 288 nsew signal input
rlabel metal2 s 78954 0 79010 800 6 wbs_adr_i[15]
port 289 nsew signal input
rlabel metal2 s 83278 0 83334 800 6 wbs_adr_i[16]
port 290 nsew signal input
rlabel metal2 s 87510 0 87566 800 6 wbs_adr_i[17]
port 291 nsew signal input
rlabel metal2 s 91834 0 91890 800 6 wbs_adr_i[18]
port 292 nsew signal input
rlabel metal2 s 96066 0 96122 800 6 wbs_adr_i[19]
port 293 nsew signal input
rlabel metal2 s 14830 0 14886 800 6 wbs_adr_i[1]
port 294 nsew signal input
rlabel metal2 s 100390 0 100446 800 6 wbs_adr_i[20]
port 295 nsew signal input
rlabel metal2 s 104622 0 104678 800 6 wbs_adr_i[21]
port 296 nsew signal input
rlabel metal2 s 108854 0 108910 800 6 wbs_adr_i[22]
port 297 nsew signal input
rlabel metal2 s 113178 0 113234 800 6 wbs_adr_i[23]
port 298 nsew signal input
rlabel metal2 s 117410 0 117466 800 6 wbs_adr_i[24]
port 299 nsew signal input
rlabel metal2 s 121734 0 121790 800 6 wbs_adr_i[25]
port 300 nsew signal input
rlabel metal2 s 125966 0 126022 800 6 wbs_adr_i[26]
port 301 nsew signal input
rlabel metal2 s 130290 0 130346 800 6 wbs_adr_i[27]
port 302 nsew signal input
rlabel metal2 s 134522 0 134578 800 6 wbs_adr_i[28]
port 303 nsew signal input
rlabel metal2 s 138846 0 138902 800 6 wbs_adr_i[29]
port 304 nsew signal input
rlabel metal2 s 20534 0 20590 800 6 wbs_adr_i[2]
port 305 nsew signal input
rlabel metal2 s 143078 0 143134 800 6 wbs_adr_i[30]
port 306 nsew signal input
rlabel metal2 s 147402 0 147458 800 6 wbs_adr_i[31]
port 307 nsew signal input
rlabel metal2 s 26238 0 26294 800 6 wbs_adr_i[3]
port 308 nsew signal input
rlabel metal2 s 31942 0 31998 800 6 wbs_adr_i[4]
port 309 nsew signal input
rlabel metal2 s 36266 0 36322 800 6 wbs_adr_i[5]
port 310 nsew signal input
rlabel metal2 s 40498 0 40554 800 6 wbs_adr_i[6]
port 311 nsew signal input
rlabel metal2 s 44822 0 44878 800 6 wbs_adr_i[7]
port 312 nsew signal input
rlabel metal2 s 49054 0 49110 800 6 wbs_adr_i[8]
port 313 nsew signal input
rlabel metal2 s 53286 0 53342 800 6 wbs_adr_i[9]
port 314 nsew signal input
rlabel metal2 s 4894 0 4950 800 6 wbs_cyc_i
port 315 nsew signal input
rlabel metal2 s 10598 0 10654 800 6 wbs_dat_i[0]
port 316 nsew signal input
rlabel metal2 s 58990 0 59046 800 6 wbs_dat_i[10]
port 317 nsew signal input
rlabel metal2 s 63314 0 63370 800 6 wbs_dat_i[11]
port 318 nsew signal input
rlabel metal2 s 67546 0 67602 800 6 wbs_dat_i[12]
port 319 nsew signal input
rlabel metal2 s 71870 0 71926 800 6 wbs_dat_i[13]
port 320 nsew signal input
rlabel metal2 s 76102 0 76158 800 6 wbs_dat_i[14]
port 321 nsew signal input
rlabel metal2 s 80426 0 80482 800 6 wbs_dat_i[15]
port 322 nsew signal input
rlabel metal2 s 84658 0 84714 800 6 wbs_dat_i[16]
port 323 nsew signal input
rlabel metal2 s 88982 0 89038 800 6 wbs_dat_i[17]
port 324 nsew signal input
rlabel metal2 s 93214 0 93270 800 6 wbs_dat_i[18]
port 325 nsew signal input
rlabel metal2 s 97538 0 97594 800 6 wbs_dat_i[19]
port 326 nsew signal input
rlabel metal2 s 16302 0 16358 800 6 wbs_dat_i[1]
port 327 nsew signal input
rlabel metal2 s 101770 0 101826 800 6 wbs_dat_i[20]
port 328 nsew signal input
rlabel metal2 s 106002 0 106058 800 6 wbs_dat_i[21]
port 329 nsew signal input
rlabel metal2 s 110326 0 110382 800 6 wbs_dat_i[22]
port 330 nsew signal input
rlabel metal2 s 114558 0 114614 800 6 wbs_dat_i[23]
port 331 nsew signal input
rlabel metal2 s 118882 0 118938 800 6 wbs_dat_i[24]
port 332 nsew signal input
rlabel metal2 s 123114 0 123170 800 6 wbs_dat_i[25]
port 333 nsew signal input
rlabel metal2 s 127438 0 127494 800 6 wbs_dat_i[26]
port 334 nsew signal input
rlabel metal2 s 131670 0 131726 800 6 wbs_dat_i[27]
port 335 nsew signal input
rlabel metal2 s 135994 0 136050 800 6 wbs_dat_i[28]
port 336 nsew signal input
rlabel metal2 s 140226 0 140282 800 6 wbs_dat_i[29]
port 337 nsew signal input
rlabel metal2 s 22006 0 22062 800 6 wbs_dat_i[2]
port 338 nsew signal input
rlabel metal2 s 144550 0 144606 800 6 wbs_dat_i[30]
port 339 nsew signal input
rlabel metal2 s 148782 0 148838 800 6 wbs_dat_i[31]
port 340 nsew signal input
rlabel metal2 s 27710 0 27766 800 6 wbs_dat_i[3]
port 341 nsew signal input
rlabel metal2 s 33414 0 33470 800 6 wbs_dat_i[4]
port 342 nsew signal input
rlabel metal2 s 37646 0 37702 800 6 wbs_dat_i[5]
port 343 nsew signal input
rlabel metal2 s 41970 0 42026 800 6 wbs_dat_i[6]
port 344 nsew signal input
rlabel metal2 s 46202 0 46258 800 6 wbs_dat_i[7]
port 345 nsew signal input
rlabel metal2 s 50526 0 50582 800 6 wbs_dat_i[8]
port 346 nsew signal input
rlabel metal2 s 54758 0 54814 800 6 wbs_dat_i[9]
port 347 nsew signal input
rlabel metal2 s 11978 0 12034 800 6 wbs_dat_o[0]
port 348 nsew signal output
rlabel metal2 s 60462 0 60518 800 6 wbs_dat_o[10]
port 349 nsew signal output
rlabel metal2 s 64694 0 64750 800 6 wbs_dat_o[11]
port 350 nsew signal output
rlabel metal2 s 69018 0 69074 800 6 wbs_dat_o[12]
port 351 nsew signal output
rlabel metal2 s 73250 0 73306 800 6 wbs_dat_o[13]
port 352 nsew signal output
rlabel metal2 s 77574 0 77630 800 6 wbs_dat_o[14]
port 353 nsew signal output
rlabel metal2 s 81806 0 81862 800 6 wbs_dat_o[15]
port 354 nsew signal output
rlabel metal2 s 86130 0 86186 800 6 wbs_dat_o[16]
port 355 nsew signal output
rlabel metal2 s 90362 0 90418 800 6 wbs_dat_o[17]
port 356 nsew signal output
rlabel metal2 s 94686 0 94742 800 6 wbs_dat_o[18]
port 357 nsew signal output
rlabel metal2 s 98918 0 98974 800 6 wbs_dat_o[19]
port 358 nsew signal output
rlabel metal2 s 17682 0 17738 800 6 wbs_dat_o[1]
port 359 nsew signal output
rlabel metal2 s 103150 0 103206 800 6 wbs_dat_o[20]
port 360 nsew signal output
rlabel metal2 s 107474 0 107530 800 6 wbs_dat_o[21]
port 361 nsew signal output
rlabel metal2 s 111706 0 111762 800 6 wbs_dat_o[22]
port 362 nsew signal output
rlabel metal2 s 116030 0 116086 800 6 wbs_dat_o[23]
port 363 nsew signal output
rlabel metal2 s 120262 0 120318 800 6 wbs_dat_o[24]
port 364 nsew signal output
rlabel metal2 s 124586 0 124642 800 6 wbs_dat_o[25]
port 365 nsew signal output
rlabel metal2 s 128818 0 128874 800 6 wbs_dat_o[26]
port 366 nsew signal output
rlabel metal2 s 133142 0 133198 800 6 wbs_dat_o[27]
port 367 nsew signal output
rlabel metal2 s 137374 0 137430 800 6 wbs_dat_o[28]
port 368 nsew signal output
rlabel metal2 s 141698 0 141754 800 6 wbs_dat_o[29]
port 369 nsew signal output
rlabel metal2 s 23386 0 23442 800 6 wbs_dat_o[2]
port 370 nsew signal output
rlabel metal2 s 145930 0 145986 800 6 wbs_dat_o[30]
port 371 nsew signal output
rlabel metal2 s 150254 0 150310 800 6 wbs_dat_o[31]
port 372 nsew signal output
rlabel metal2 s 29090 0 29146 800 6 wbs_dat_o[3]
port 373 nsew signal output
rlabel metal2 s 34794 0 34850 800 6 wbs_dat_o[4]
port 374 nsew signal output
rlabel metal2 s 39118 0 39174 800 6 wbs_dat_o[5]
port 375 nsew signal output
rlabel metal2 s 43350 0 43406 800 6 wbs_dat_o[6]
port 376 nsew signal output
rlabel metal2 s 47674 0 47730 800 6 wbs_dat_o[7]
port 377 nsew signal output
rlabel metal2 s 51906 0 51962 800 6 wbs_dat_o[8]
port 378 nsew signal output
rlabel metal2 s 56138 0 56194 800 6 wbs_dat_o[9]
port 379 nsew signal output
rlabel metal2 s 13450 0 13506 800 6 wbs_sel_i[0]
port 380 nsew signal input
rlabel metal2 s 19154 0 19210 800 6 wbs_sel_i[1]
port 381 nsew signal input
rlabel metal2 s 24858 0 24914 800 6 wbs_sel_i[2]
port 382 nsew signal input
rlabel metal2 s 30562 0 30618 800 6 wbs_sel_i[3]
port 383 nsew signal input
rlabel metal2 s 6274 0 6330 800 6 wbs_stb_i
port 384 nsew signal input
rlabel metal2 s 7746 0 7802 800 6 wbs_we_i
port 385 nsew signal input
<< properties >>
string LEFclass BLOCK
string FIXED_BBOX 0 0 199424 201568
string LEFview TRUE
string GDS_FILE /local/home/roman/projects/opencircuitdesign/shuttle5/caravel_mpw/openlane/user_proj/runs/user_proj/results/magic/user_proj.gds
string GDS_END 99314092
string GDS_START 1436846
<< end >>

