magic
tech sky130A
magscale 1 2
timestamp 1641262152
<< obsli1 >>
rect 1104 1445 178451 180523
<< obsm1 >>
rect 566 756 178650 180792
<< metal2 >>
rect 570 180003 626 180803
rect 1674 180003 1730 180803
rect 2870 180003 2926 180803
rect 4066 180003 4122 180803
rect 5262 180003 5318 180803
rect 6458 180003 6514 180803
rect 7654 180003 7710 180803
rect 8850 180003 8906 180803
rect 10046 180003 10102 180803
rect 11242 180003 11298 180803
rect 12438 180003 12494 180803
rect 13634 180003 13690 180803
rect 14830 180003 14886 180803
rect 16026 180003 16082 180803
rect 17222 180003 17278 180803
rect 18418 180003 18474 180803
rect 19614 180003 19670 180803
rect 20810 180003 20866 180803
rect 22006 180003 22062 180803
rect 23110 180003 23166 180803
rect 24306 180003 24362 180803
rect 25502 180003 25558 180803
rect 26698 180003 26754 180803
rect 27894 180003 27950 180803
rect 29090 180003 29146 180803
rect 30286 180003 30342 180803
rect 31482 180003 31538 180803
rect 32678 180003 32734 180803
rect 33874 180003 33930 180803
rect 35070 180003 35126 180803
rect 36266 180003 36322 180803
rect 37462 180003 37518 180803
rect 38658 180003 38714 180803
rect 39854 180003 39910 180803
rect 41050 180003 41106 180803
rect 42246 180003 42302 180803
rect 43442 180003 43498 180803
rect 44638 180003 44694 180803
rect 45742 180003 45798 180803
rect 46938 180003 46994 180803
rect 48134 180003 48190 180803
rect 49330 180003 49386 180803
rect 50526 180003 50582 180803
rect 51722 180003 51778 180803
rect 52918 180003 52974 180803
rect 54114 180003 54170 180803
rect 55310 180003 55366 180803
rect 56506 180003 56562 180803
rect 57702 180003 57758 180803
rect 58898 180003 58954 180803
rect 60094 180003 60150 180803
rect 61290 180003 61346 180803
rect 62486 180003 62542 180803
rect 63682 180003 63738 180803
rect 64878 180003 64934 180803
rect 66074 180003 66130 180803
rect 67270 180003 67326 180803
rect 68374 180003 68430 180803
rect 69570 180003 69626 180803
rect 70766 180003 70822 180803
rect 71962 180003 72018 180803
rect 73158 180003 73214 180803
rect 74354 180003 74410 180803
rect 75550 180003 75606 180803
rect 76746 180003 76802 180803
rect 77942 180003 77998 180803
rect 79138 180003 79194 180803
rect 80334 180003 80390 180803
rect 81530 180003 81586 180803
rect 82726 180003 82782 180803
rect 83922 180003 83978 180803
rect 85118 180003 85174 180803
rect 86314 180003 86370 180803
rect 87510 180003 87566 180803
rect 88706 180003 88762 180803
rect 89902 180003 89958 180803
rect 91006 180003 91062 180803
rect 92202 180003 92258 180803
rect 93398 180003 93454 180803
rect 94594 180003 94650 180803
rect 95790 180003 95846 180803
rect 96986 180003 97042 180803
rect 98182 180003 98238 180803
rect 99378 180003 99434 180803
rect 100574 180003 100630 180803
rect 101770 180003 101826 180803
rect 102966 180003 103022 180803
rect 104162 180003 104218 180803
rect 105358 180003 105414 180803
rect 106554 180003 106610 180803
rect 107750 180003 107806 180803
rect 108946 180003 109002 180803
rect 110142 180003 110198 180803
rect 111338 180003 111394 180803
rect 112442 180003 112498 180803
rect 113638 180003 113694 180803
rect 114834 180003 114890 180803
rect 116030 180003 116086 180803
rect 117226 180003 117282 180803
rect 118422 180003 118478 180803
rect 119618 180003 119674 180803
rect 120814 180003 120870 180803
rect 122010 180003 122066 180803
rect 123206 180003 123262 180803
rect 124402 180003 124458 180803
rect 125598 180003 125654 180803
rect 126794 180003 126850 180803
rect 127990 180003 128046 180803
rect 129186 180003 129242 180803
rect 130382 180003 130438 180803
rect 131578 180003 131634 180803
rect 132774 180003 132830 180803
rect 133970 180003 134026 180803
rect 135074 180003 135130 180803
rect 136270 180003 136326 180803
rect 137466 180003 137522 180803
rect 138662 180003 138718 180803
rect 139858 180003 139914 180803
rect 141054 180003 141110 180803
rect 142250 180003 142306 180803
rect 143446 180003 143502 180803
rect 144642 180003 144698 180803
rect 145838 180003 145894 180803
rect 147034 180003 147090 180803
rect 148230 180003 148286 180803
rect 149426 180003 149482 180803
rect 150622 180003 150678 180803
rect 151818 180003 151874 180803
rect 153014 180003 153070 180803
rect 154210 180003 154266 180803
rect 155406 180003 155462 180803
rect 156602 180003 156658 180803
rect 157706 180003 157762 180803
rect 158902 180003 158958 180803
rect 160098 180003 160154 180803
rect 161294 180003 161350 180803
rect 162490 180003 162546 180803
rect 163686 180003 163742 180803
rect 164882 180003 164938 180803
rect 166078 180003 166134 180803
rect 167274 180003 167330 180803
rect 168470 180003 168526 180803
rect 169666 180003 169722 180803
rect 170862 180003 170918 180803
rect 172058 180003 172114 180803
rect 173254 180003 173310 180803
rect 174450 180003 174506 180803
rect 175646 180003 175702 180803
rect 176842 180003 176898 180803
rect 178038 180003 178094 180803
rect 570 0 626 800
rect 1766 0 1822 800
rect 2962 0 3018 800
rect 4158 0 4214 800
rect 5446 0 5502 800
rect 6642 0 6698 800
rect 7838 0 7894 800
rect 9126 0 9182 800
rect 10322 0 10378 800
rect 11518 0 11574 800
rect 12806 0 12862 800
rect 14002 0 14058 800
rect 15198 0 15254 800
rect 16394 0 16450 800
rect 17682 0 17738 800
rect 18878 0 18934 800
rect 20074 0 20130 800
rect 21362 0 21418 800
rect 22558 0 22614 800
rect 23754 0 23810 800
rect 25042 0 25098 800
rect 26238 0 26294 800
rect 27434 0 27490 800
rect 28630 0 28686 800
rect 29918 0 29974 800
rect 31114 0 31170 800
rect 32310 0 32366 800
rect 33598 0 33654 800
rect 34794 0 34850 800
rect 35990 0 36046 800
rect 37278 0 37334 800
rect 38474 0 38530 800
rect 39670 0 39726 800
rect 40866 0 40922 800
rect 42154 0 42210 800
rect 43350 0 43406 800
rect 44546 0 44602 800
rect 45834 0 45890 800
rect 47030 0 47086 800
rect 48226 0 48282 800
rect 49514 0 49570 800
rect 50710 0 50766 800
rect 51906 0 51962 800
rect 53102 0 53158 800
rect 54390 0 54446 800
rect 55586 0 55642 800
rect 56782 0 56838 800
rect 58070 0 58126 800
rect 59266 0 59322 800
rect 60462 0 60518 800
rect 61750 0 61806 800
rect 62946 0 63002 800
rect 64142 0 64198 800
rect 65338 0 65394 800
rect 66626 0 66682 800
rect 67822 0 67878 800
rect 69018 0 69074 800
rect 70306 0 70362 800
rect 71502 0 71558 800
rect 72698 0 72754 800
rect 73986 0 74042 800
rect 75182 0 75238 800
rect 76378 0 76434 800
rect 77574 0 77630 800
rect 78862 0 78918 800
rect 80058 0 80114 800
rect 81254 0 81310 800
rect 82542 0 82598 800
rect 83738 0 83794 800
rect 84934 0 84990 800
rect 86222 0 86278 800
rect 87418 0 87474 800
rect 88614 0 88670 800
rect 89902 0 89958 800
rect 91098 0 91154 800
rect 92294 0 92350 800
rect 93490 0 93546 800
rect 94778 0 94834 800
rect 95974 0 96030 800
rect 97170 0 97226 800
rect 98458 0 98514 800
rect 99654 0 99710 800
rect 100850 0 100906 800
rect 102138 0 102194 800
rect 103334 0 103390 800
rect 104530 0 104586 800
rect 105726 0 105782 800
rect 107014 0 107070 800
rect 108210 0 108266 800
rect 109406 0 109462 800
rect 110694 0 110750 800
rect 111890 0 111946 800
rect 113086 0 113142 800
rect 114374 0 114430 800
rect 115570 0 115626 800
rect 116766 0 116822 800
rect 117962 0 118018 800
rect 119250 0 119306 800
rect 120446 0 120502 800
rect 121642 0 121698 800
rect 122930 0 122986 800
rect 124126 0 124182 800
rect 125322 0 125378 800
rect 126610 0 126666 800
rect 127806 0 127862 800
rect 129002 0 129058 800
rect 130198 0 130254 800
rect 131486 0 131542 800
rect 132682 0 132738 800
rect 133878 0 133934 800
rect 135166 0 135222 800
rect 136362 0 136418 800
rect 137558 0 137614 800
rect 138846 0 138902 800
rect 140042 0 140098 800
rect 141238 0 141294 800
rect 142434 0 142490 800
rect 143722 0 143778 800
rect 144918 0 144974 800
rect 146114 0 146170 800
rect 147402 0 147458 800
rect 148598 0 148654 800
rect 149794 0 149850 800
rect 151082 0 151138 800
rect 152278 0 152334 800
rect 153474 0 153530 800
rect 154670 0 154726 800
rect 155958 0 156014 800
rect 157154 0 157210 800
rect 158350 0 158406 800
rect 159638 0 159694 800
rect 160834 0 160890 800
rect 162030 0 162086 800
rect 163318 0 163374 800
rect 164514 0 164570 800
rect 165710 0 165766 800
rect 166906 0 166962 800
rect 168194 0 168250 800
rect 169390 0 169446 800
rect 170586 0 170642 800
rect 171874 0 171930 800
rect 173070 0 173126 800
rect 174266 0 174322 800
rect 175554 0 175610 800
rect 176750 0 176806 800
rect 177946 0 178002 800
<< obsm2 >>
rect 682 179947 1618 180742
rect 1786 179947 2814 180742
rect 2982 179947 4010 180742
rect 4178 179947 5206 180742
rect 5374 179947 6402 180742
rect 6570 179947 7598 180742
rect 7766 179947 8794 180742
rect 8962 179947 9990 180742
rect 10158 179947 11186 180742
rect 11354 179947 12382 180742
rect 12550 179947 13578 180742
rect 13746 179947 14774 180742
rect 14942 179947 15970 180742
rect 16138 179947 17166 180742
rect 17334 179947 18362 180742
rect 18530 179947 19558 180742
rect 19726 179947 20754 180742
rect 20922 179947 21950 180742
rect 22118 179947 23054 180742
rect 23222 179947 24250 180742
rect 24418 179947 25446 180742
rect 25614 179947 26642 180742
rect 26810 179947 27838 180742
rect 28006 179947 29034 180742
rect 29202 179947 30230 180742
rect 30398 179947 31426 180742
rect 31594 179947 32622 180742
rect 32790 179947 33818 180742
rect 33986 179947 35014 180742
rect 35182 179947 36210 180742
rect 36378 179947 37406 180742
rect 37574 179947 38602 180742
rect 38770 179947 39798 180742
rect 39966 179947 40994 180742
rect 41162 179947 42190 180742
rect 42358 179947 43386 180742
rect 43554 179947 44582 180742
rect 44750 179947 45686 180742
rect 45854 179947 46882 180742
rect 47050 179947 48078 180742
rect 48246 179947 49274 180742
rect 49442 179947 50470 180742
rect 50638 179947 51666 180742
rect 51834 179947 52862 180742
rect 53030 179947 54058 180742
rect 54226 179947 55254 180742
rect 55422 179947 56450 180742
rect 56618 179947 57646 180742
rect 57814 179947 58842 180742
rect 59010 179947 60038 180742
rect 60206 179947 61234 180742
rect 61402 179947 62430 180742
rect 62598 179947 63626 180742
rect 63794 179947 64822 180742
rect 64990 179947 66018 180742
rect 66186 179947 67214 180742
rect 67382 179947 68318 180742
rect 68486 179947 69514 180742
rect 69682 179947 70710 180742
rect 70878 179947 71906 180742
rect 72074 179947 73102 180742
rect 73270 179947 74298 180742
rect 74466 179947 75494 180742
rect 75662 179947 76690 180742
rect 76858 179947 77886 180742
rect 78054 179947 79082 180742
rect 79250 179947 80278 180742
rect 80446 179947 81474 180742
rect 81642 179947 82670 180742
rect 82838 179947 83866 180742
rect 84034 179947 85062 180742
rect 85230 179947 86258 180742
rect 86426 179947 87454 180742
rect 87622 179947 88650 180742
rect 88818 179947 89846 180742
rect 90014 179947 90950 180742
rect 91118 179947 92146 180742
rect 92314 179947 93342 180742
rect 93510 179947 94538 180742
rect 94706 179947 95734 180742
rect 95902 179947 96930 180742
rect 97098 179947 98126 180742
rect 98294 179947 99322 180742
rect 99490 179947 100518 180742
rect 100686 179947 101714 180742
rect 101882 179947 102910 180742
rect 103078 179947 104106 180742
rect 104274 179947 105302 180742
rect 105470 179947 106498 180742
rect 106666 179947 107694 180742
rect 107862 179947 108890 180742
rect 109058 179947 110086 180742
rect 110254 179947 111282 180742
rect 111450 179947 112386 180742
rect 112554 179947 113582 180742
rect 113750 179947 114778 180742
rect 114946 179947 115974 180742
rect 116142 179947 117170 180742
rect 117338 179947 118366 180742
rect 118534 179947 119562 180742
rect 119730 179947 120758 180742
rect 120926 179947 121954 180742
rect 122122 179947 123150 180742
rect 123318 179947 124346 180742
rect 124514 179947 125542 180742
rect 125710 179947 126738 180742
rect 126906 179947 127934 180742
rect 128102 179947 129130 180742
rect 129298 179947 130326 180742
rect 130494 179947 131522 180742
rect 131690 179947 132718 180742
rect 132886 179947 133914 180742
rect 134082 179947 135018 180742
rect 135186 179947 136214 180742
rect 136382 179947 137410 180742
rect 137578 179947 138606 180742
rect 138774 179947 139802 180742
rect 139970 179947 140998 180742
rect 141166 179947 142194 180742
rect 142362 179947 143390 180742
rect 143558 179947 144586 180742
rect 144754 179947 145782 180742
rect 145950 179947 146978 180742
rect 147146 179947 148174 180742
rect 148342 179947 149370 180742
rect 149538 179947 150566 180742
rect 150734 179947 151762 180742
rect 151930 179947 152958 180742
rect 153126 179947 154154 180742
rect 154322 179947 155350 180742
rect 155518 179947 156546 180742
rect 156714 179947 157650 180742
rect 157818 179947 158846 180742
rect 159014 179947 160042 180742
rect 160210 179947 161238 180742
rect 161406 179947 162434 180742
rect 162602 179947 163630 180742
rect 163798 179947 164826 180742
rect 164994 179947 166022 180742
rect 166190 179947 167218 180742
rect 167386 179947 168414 180742
rect 168582 179947 169610 180742
rect 169778 179947 170806 180742
rect 170974 179947 172002 180742
rect 172170 179947 173198 180742
rect 173366 179947 174394 180742
rect 174562 179947 175590 180742
rect 175758 179947 176786 180742
rect 176954 179947 177982 180742
rect 178150 179947 178646 180742
rect 572 856 178646 179947
rect 682 734 1710 856
rect 1878 734 2906 856
rect 3074 734 4102 856
rect 4270 734 5390 856
rect 5558 734 6586 856
rect 6754 734 7782 856
rect 7950 734 9070 856
rect 9238 734 10266 856
rect 10434 734 11462 856
rect 11630 734 12750 856
rect 12918 734 13946 856
rect 14114 734 15142 856
rect 15310 734 16338 856
rect 16506 734 17626 856
rect 17794 734 18822 856
rect 18990 734 20018 856
rect 20186 734 21306 856
rect 21474 734 22502 856
rect 22670 734 23698 856
rect 23866 734 24986 856
rect 25154 734 26182 856
rect 26350 734 27378 856
rect 27546 734 28574 856
rect 28742 734 29862 856
rect 30030 734 31058 856
rect 31226 734 32254 856
rect 32422 734 33542 856
rect 33710 734 34738 856
rect 34906 734 35934 856
rect 36102 734 37222 856
rect 37390 734 38418 856
rect 38586 734 39614 856
rect 39782 734 40810 856
rect 40978 734 42098 856
rect 42266 734 43294 856
rect 43462 734 44490 856
rect 44658 734 45778 856
rect 45946 734 46974 856
rect 47142 734 48170 856
rect 48338 734 49458 856
rect 49626 734 50654 856
rect 50822 734 51850 856
rect 52018 734 53046 856
rect 53214 734 54334 856
rect 54502 734 55530 856
rect 55698 734 56726 856
rect 56894 734 58014 856
rect 58182 734 59210 856
rect 59378 734 60406 856
rect 60574 734 61694 856
rect 61862 734 62890 856
rect 63058 734 64086 856
rect 64254 734 65282 856
rect 65450 734 66570 856
rect 66738 734 67766 856
rect 67934 734 68962 856
rect 69130 734 70250 856
rect 70418 734 71446 856
rect 71614 734 72642 856
rect 72810 734 73930 856
rect 74098 734 75126 856
rect 75294 734 76322 856
rect 76490 734 77518 856
rect 77686 734 78806 856
rect 78974 734 80002 856
rect 80170 734 81198 856
rect 81366 734 82486 856
rect 82654 734 83682 856
rect 83850 734 84878 856
rect 85046 734 86166 856
rect 86334 734 87362 856
rect 87530 734 88558 856
rect 88726 734 89846 856
rect 90014 734 91042 856
rect 91210 734 92238 856
rect 92406 734 93434 856
rect 93602 734 94722 856
rect 94890 734 95918 856
rect 96086 734 97114 856
rect 97282 734 98402 856
rect 98570 734 99598 856
rect 99766 734 100794 856
rect 100962 734 102082 856
rect 102250 734 103278 856
rect 103446 734 104474 856
rect 104642 734 105670 856
rect 105838 734 106958 856
rect 107126 734 108154 856
rect 108322 734 109350 856
rect 109518 734 110638 856
rect 110806 734 111834 856
rect 112002 734 113030 856
rect 113198 734 114318 856
rect 114486 734 115514 856
rect 115682 734 116710 856
rect 116878 734 117906 856
rect 118074 734 119194 856
rect 119362 734 120390 856
rect 120558 734 121586 856
rect 121754 734 122874 856
rect 123042 734 124070 856
rect 124238 734 125266 856
rect 125434 734 126554 856
rect 126722 734 127750 856
rect 127918 734 128946 856
rect 129114 734 130142 856
rect 130310 734 131430 856
rect 131598 734 132626 856
rect 132794 734 133822 856
rect 133990 734 135110 856
rect 135278 734 136306 856
rect 136474 734 137502 856
rect 137670 734 138790 856
rect 138958 734 139986 856
rect 140154 734 141182 856
rect 141350 734 142378 856
rect 142546 734 143666 856
rect 143834 734 144862 856
rect 145030 734 146058 856
rect 146226 734 147346 856
rect 147514 734 148542 856
rect 148710 734 149738 856
rect 149906 734 151026 856
rect 151194 734 152222 856
rect 152390 734 153418 856
rect 153586 734 154614 856
rect 154782 734 155902 856
rect 156070 734 157098 856
rect 157266 734 158294 856
rect 158462 734 159582 856
rect 159750 734 160778 856
rect 160946 734 161974 856
rect 162142 734 163262 856
rect 163430 734 164458 856
rect 164626 734 165654 856
rect 165822 734 166850 856
rect 167018 734 168138 856
rect 168306 734 169334 856
rect 169502 734 170530 856
rect 170698 734 171818 856
rect 171986 734 173014 856
rect 173182 734 174210 856
rect 174378 734 175498 856
rect 175666 734 176694 856
rect 176862 734 177890 856
rect 178058 734 178646 856
<< metal3 >>
rect 177859 178712 178659 178832
rect 0 178440 800 178560
rect 177859 174768 178659 174888
rect 0 174088 800 174208
rect 177859 170824 178659 170944
rect 0 169600 800 169720
rect 177859 166880 178659 167000
rect 0 165248 800 165368
rect 177859 162936 178659 163056
rect 0 160760 800 160880
rect 177859 158992 178659 159112
rect 0 156408 800 156528
rect 177859 155048 178659 155168
rect 0 152056 800 152176
rect 177859 151104 178659 151224
rect 0 147568 800 147688
rect 177859 147160 178659 147280
rect 0 143216 800 143336
rect 177859 143352 178659 143472
rect 177859 139408 178659 139528
rect 0 138728 800 138848
rect 177859 135464 178659 135584
rect 0 134376 800 134496
rect 177859 131520 178659 131640
rect 0 130024 800 130144
rect 177859 127576 178659 127696
rect 0 125536 800 125656
rect 177859 123632 178659 123752
rect 0 121184 800 121304
rect 177859 119688 178659 119808
rect 0 116696 800 116816
rect 177859 115744 178659 115864
rect 0 112344 800 112464
rect 177859 111800 178659 111920
rect 0 107856 800 107976
rect 177859 107992 178659 108112
rect 177859 104048 178659 104168
rect 0 103504 800 103624
rect 177859 100104 178659 100224
rect 0 99152 800 99272
rect 177859 96160 178659 96280
rect 0 94664 800 94784
rect 177859 92216 178659 92336
rect 0 90312 800 90432
rect 177859 88272 178659 88392
rect 0 85824 800 85944
rect 177859 84328 178659 84448
rect 0 81472 800 81592
rect 177859 80384 178659 80504
rect 0 77120 800 77240
rect 177859 76440 178659 76560
rect 0 72632 800 72752
rect 177859 72632 178659 72752
rect 177859 68688 178659 68808
rect 0 68280 800 68400
rect 177859 64744 178659 64864
rect 0 63792 800 63912
rect 177859 60800 178659 60920
rect 0 59440 800 59560
rect 177859 56856 178659 56976
rect 0 54952 800 55072
rect 177859 52912 178659 53032
rect 0 50600 800 50720
rect 177859 48968 178659 49088
rect 0 46248 800 46368
rect 177859 45024 178659 45144
rect 0 41760 800 41880
rect 177859 41080 178659 41200
rect 0 37408 800 37528
rect 177859 37272 178659 37392
rect 177859 33328 178659 33448
rect 0 32920 800 33040
rect 177859 29384 178659 29504
rect 0 28568 800 28688
rect 177859 25440 178659 25560
rect 0 24216 800 24336
rect 177859 21496 178659 21616
rect 0 19728 800 19848
rect 177859 17552 178659 17672
rect 0 15376 800 15496
rect 177859 13608 178659 13728
rect 0 10888 800 11008
rect 177859 9664 178659 9784
rect 0 6536 800 6656
rect 177859 5720 178659 5840
rect 0 2184 800 2304
rect 177859 1912 178659 2032
<< obsm3 >>
rect 800 178912 178651 180709
rect 800 178640 177779 178912
rect 880 178632 177779 178640
rect 880 178360 178651 178632
rect 800 174968 178651 178360
rect 800 174688 177779 174968
rect 800 174288 178651 174688
rect 880 174008 178651 174288
rect 800 171024 178651 174008
rect 800 170744 177779 171024
rect 800 169800 178651 170744
rect 880 169520 178651 169800
rect 800 167080 178651 169520
rect 800 166800 177779 167080
rect 800 165448 178651 166800
rect 880 165168 178651 165448
rect 800 163136 178651 165168
rect 800 162856 177779 163136
rect 800 160960 178651 162856
rect 880 160680 178651 160960
rect 800 159192 178651 160680
rect 800 158912 177779 159192
rect 800 156608 178651 158912
rect 880 156328 178651 156608
rect 800 155248 178651 156328
rect 800 154968 177779 155248
rect 800 152256 178651 154968
rect 880 151976 178651 152256
rect 800 151304 178651 151976
rect 800 151024 177779 151304
rect 800 147768 178651 151024
rect 880 147488 178651 147768
rect 800 147360 178651 147488
rect 800 147080 177779 147360
rect 800 143552 178651 147080
rect 800 143416 177779 143552
rect 880 143272 177779 143416
rect 880 143136 178651 143272
rect 800 139608 178651 143136
rect 800 139328 177779 139608
rect 800 138928 178651 139328
rect 880 138648 178651 138928
rect 800 135664 178651 138648
rect 800 135384 177779 135664
rect 800 134576 178651 135384
rect 880 134296 178651 134576
rect 800 131720 178651 134296
rect 800 131440 177779 131720
rect 800 130224 178651 131440
rect 880 129944 178651 130224
rect 800 127776 178651 129944
rect 800 127496 177779 127776
rect 800 125736 178651 127496
rect 880 125456 178651 125736
rect 800 123832 178651 125456
rect 800 123552 177779 123832
rect 800 121384 178651 123552
rect 880 121104 178651 121384
rect 800 119888 178651 121104
rect 800 119608 177779 119888
rect 800 116896 178651 119608
rect 880 116616 178651 116896
rect 800 115944 178651 116616
rect 800 115664 177779 115944
rect 800 112544 178651 115664
rect 880 112264 178651 112544
rect 800 112000 178651 112264
rect 800 111720 177779 112000
rect 800 108192 178651 111720
rect 800 108056 177779 108192
rect 880 107912 177779 108056
rect 880 107776 178651 107912
rect 800 104248 178651 107776
rect 800 103968 177779 104248
rect 800 103704 178651 103968
rect 880 103424 178651 103704
rect 800 100304 178651 103424
rect 800 100024 177779 100304
rect 800 99352 178651 100024
rect 880 99072 178651 99352
rect 800 96360 178651 99072
rect 800 96080 177779 96360
rect 800 94864 178651 96080
rect 880 94584 178651 94864
rect 800 92416 178651 94584
rect 800 92136 177779 92416
rect 800 90512 178651 92136
rect 880 90232 178651 90512
rect 800 88472 178651 90232
rect 800 88192 177779 88472
rect 800 86024 178651 88192
rect 880 85744 178651 86024
rect 800 84528 178651 85744
rect 800 84248 177779 84528
rect 800 81672 178651 84248
rect 880 81392 178651 81672
rect 800 80584 178651 81392
rect 800 80304 177779 80584
rect 800 77320 178651 80304
rect 880 77040 178651 77320
rect 800 76640 178651 77040
rect 800 76360 177779 76640
rect 800 72832 178651 76360
rect 880 72552 177779 72832
rect 800 68888 178651 72552
rect 800 68608 177779 68888
rect 800 68480 178651 68608
rect 880 68200 178651 68480
rect 800 64944 178651 68200
rect 800 64664 177779 64944
rect 800 63992 178651 64664
rect 880 63712 178651 63992
rect 800 61000 178651 63712
rect 800 60720 177779 61000
rect 800 59640 178651 60720
rect 880 59360 178651 59640
rect 800 57056 178651 59360
rect 800 56776 177779 57056
rect 800 55152 178651 56776
rect 880 54872 178651 55152
rect 800 53112 178651 54872
rect 800 52832 177779 53112
rect 800 50800 178651 52832
rect 880 50520 178651 50800
rect 800 49168 178651 50520
rect 800 48888 177779 49168
rect 800 46448 178651 48888
rect 880 46168 178651 46448
rect 800 45224 178651 46168
rect 800 44944 177779 45224
rect 800 41960 178651 44944
rect 880 41680 178651 41960
rect 800 41280 178651 41680
rect 800 41000 177779 41280
rect 800 37608 178651 41000
rect 880 37472 178651 37608
rect 880 37328 177779 37472
rect 800 37192 177779 37328
rect 800 33528 178651 37192
rect 800 33248 177779 33528
rect 800 33120 178651 33248
rect 880 32840 178651 33120
rect 800 29584 178651 32840
rect 800 29304 177779 29584
rect 800 28768 178651 29304
rect 880 28488 178651 28768
rect 800 25640 178651 28488
rect 800 25360 177779 25640
rect 800 24416 178651 25360
rect 880 24136 178651 24416
rect 800 21696 178651 24136
rect 800 21416 177779 21696
rect 800 19928 178651 21416
rect 880 19648 178651 19928
rect 800 17752 178651 19648
rect 800 17472 177779 17752
rect 800 15576 178651 17472
rect 880 15296 178651 15576
rect 800 13808 178651 15296
rect 800 13528 177779 13808
rect 800 11088 178651 13528
rect 880 10808 178651 11088
rect 800 9864 178651 10808
rect 800 9584 177779 9864
rect 800 6736 178651 9584
rect 880 6456 178651 6736
rect 800 5920 178651 6456
rect 800 5640 177779 5920
rect 800 2384 178651 5640
rect 880 2112 178651 2384
rect 880 2104 177779 2112
rect 800 1832 177779 2104
rect 800 1803 178651 1832
<< metal4 >>
rect 4208 2128 4528 178480
rect 19568 2128 19888 178480
rect 34928 2128 35248 178480
rect 50288 2128 50608 178480
rect 65648 2128 65968 178480
rect 81008 2128 81328 178480
rect 96368 2128 96688 178480
rect 111728 2128 112048 178480
rect 127088 2128 127408 178480
rect 142448 2128 142768 178480
rect 157808 2128 158128 178480
rect 173168 2128 173488 178480
<< obsm4 >>
rect 6131 178560 176213 180709
rect 6131 4795 19488 178560
rect 19968 4795 34848 178560
rect 35328 4795 50208 178560
rect 50688 4795 65568 178560
rect 66048 4795 80928 178560
rect 81408 4795 96288 178560
rect 96768 4795 111648 178560
rect 112128 4795 127008 178560
rect 127488 4795 142368 178560
rect 142848 4795 157728 178560
rect 158208 4795 173088 178560
rect 173568 4795 176213 178560
<< labels >>
rlabel metal2 s 133878 0 133934 800 6 clk_i
port 1 nsew signal input
rlabel metal3 s 177859 5720 178659 5840 6 i_dout0[0]
port 2 nsew signal input
rlabel metal3 s 177859 104048 178659 104168 6 i_dout0[10]
port 3 nsew signal input
rlabel metal2 s 155958 0 156014 800 6 i_dout0[11]
port 4 nsew signal input
rlabel metal3 s 177859 111800 178659 111920 6 i_dout0[12]
port 5 nsew signal input
rlabel metal2 s 158350 0 158406 800 6 i_dout0[13]
port 6 nsew signal input
rlabel metal2 s 156602 180003 156658 180803 6 i_dout0[14]
port 7 nsew signal input
rlabel metal2 s 160834 0 160890 800 6 i_dout0[15]
port 8 nsew signal input
rlabel metal2 s 163318 0 163374 800 6 i_dout0[16]
port 9 nsew signal input
rlabel metal2 s 166906 0 166962 800 6 i_dout0[17]
port 10 nsew signal input
rlabel metal2 s 161294 180003 161350 180803 6 i_dout0[18]
port 11 nsew signal input
rlabel metal2 s 162490 180003 162546 180803 6 i_dout0[19]
port 12 nsew signal input
rlabel metal3 s 0 15376 800 15496 6 i_dout0[1]
port 13 nsew signal input
rlabel metal3 s 177859 139408 178659 139528 6 i_dout0[20]
port 14 nsew signal input
rlabel metal3 s 0 125536 800 125656 6 i_dout0[21]
port 15 nsew signal input
rlabel metal2 s 168194 0 168250 800 6 i_dout0[22]
port 16 nsew signal input
rlabel metal2 s 168470 180003 168526 180803 6 i_dout0[23]
port 17 nsew signal input
rlabel metal3 s 0 143216 800 143336 6 i_dout0[24]
port 18 nsew signal input
rlabel metal3 s 177859 158992 178659 159112 6 i_dout0[25]
port 19 nsew signal input
rlabel metal2 s 172058 180003 172114 180803 6 i_dout0[26]
port 20 nsew signal input
rlabel metal2 s 174266 0 174322 800 6 i_dout0[27]
port 21 nsew signal input
rlabel metal3 s 0 160760 800 160880 6 i_dout0[28]
port 22 nsew signal input
rlabel metal3 s 0 174088 800 174208 6 i_dout0[29]
port 23 nsew signal input
rlabel metal3 s 177859 41080 178659 41200 6 i_dout0[2]
port 24 nsew signal input
rlabel metal2 s 174450 180003 174506 180803 6 i_dout0[30]
port 25 nsew signal input
rlabel metal2 s 177946 0 178002 800 6 i_dout0[31]
port 26 nsew signal input
rlabel metal3 s 0 24216 800 24336 6 i_dout0[3]
port 27 nsew signal input
rlabel metal3 s 177859 64744 178659 64864 6 i_dout0[4]
port 28 nsew signal input
rlabel metal2 s 142434 0 142490 800 6 i_dout0[5]
port 29 nsew signal input
rlabel metal3 s 0 54952 800 55072 6 i_dout0[6]
port 30 nsew signal input
rlabel metal2 s 147034 180003 147090 180803 6 i_dout0[7]
port 31 nsew signal input
rlabel metal2 s 149794 0 149850 800 6 i_dout0[8]
port 32 nsew signal input
rlabel metal3 s 177859 100104 178659 100224 6 i_dout0[9]
port 33 nsew signal input
rlabel metal2 s 137466 180003 137522 180803 6 i_dout0_1[0]
port 34 nsew signal input
rlabel metal2 s 152278 0 152334 800 6 i_dout0_1[10]
port 35 nsew signal input
rlabel metal3 s 0 81472 800 81592 6 i_dout0_1[11]
port 36 nsew signal input
rlabel metal3 s 177859 107992 178659 108112 6 i_dout0_1[12]
port 37 nsew signal input
rlabel metal2 s 154210 180003 154266 180803 6 i_dout0_1[13]
port 38 nsew signal input
rlabel metal2 s 155406 180003 155462 180803 6 i_dout0_1[14]
port 39 nsew signal input
rlabel metal2 s 158902 180003 158958 180803 6 i_dout0_1[15]
port 40 nsew signal input
rlabel metal3 s 0 99152 800 99272 6 i_dout0_1[16]
port 41 nsew signal input
rlabel metal2 s 165710 0 165766 800 6 i_dout0_1[17]
port 42 nsew signal input
rlabel metal3 s 177859 127576 178659 127696 6 i_dout0_1[18]
port 43 nsew signal input
rlabel metal3 s 0 112344 800 112464 6 i_dout0_1[19]
port 44 nsew signal input
rlabel metal3 s 177859 25440 178659 25560 6 i_dout0_1[1]
port 45 nsew signal input
rlabel metal2 s 163686 180003 163742 180803 6 i_dout0_1[20]
port 46 nsew signal input
rlabel metal2 s 164882 180003 164938 180803 6 i_dout0_1[21]
port 47 nsew signal input
rlabel metal3 s 0 134376 800 134496 6 i_dout0_1[22]
port 48 nsew signal input
rlabel metal2 s 169390 0 169446 800 6 i_dout0_1[23]
port 49 nsew signal input
rlabel metal3 s 177859 151104 178659 151224 6 i_dout0_1[24]
port 50 nsew signal input
rlabel metal2 s 170862 180003 170918 180803 6 i_dout0_1[25]
port 51 nsew signal input
rlabel metal3 s 0 152056 800 152176 6 i_dout0_1[26]
port 52 nsew signal input
rlabel metal2 s 173070 0 173126 800 6 i_dout0_1[27]
port 53 nsew signal input
rlabel metal3 s 0 156408 800 156528 6 i_dout0_1[28]
port 54 nsew signal input
rlabel metal2 s 173254 180003 173310 180803 6 i_dout0_1[29]
port 55 nsew signal input
rlabel metal3 s 177859 37272 178659 37392 6 i_dout0_1[2]
port 56 nsew signal input
rlabel metal3 s 0 178440 800 178560 6 i_dout0_1[30]
port 57 nsew signal input
rlabel metal3 s 177859 178712 178659 178832 6 i_dout0_1[31]
port 58 nsew signal input
rlabel metal3 s 177859 48968 178659 49088 6 i_dout0_1[3]
port 59 nsew signal input
rlabel metal2 s 144642 180003 144698 180803 6 i_dout0_1[4]
port 60 nsew signal input
rlabel metal2 s 141238 0 141294 800 6 i_dout0_1[5]
port 61 nsew signal input
rlabel metal3 s 177859 76440 178659 76560 6 i_dout0_1[6]
port 62 nsew signal input
rlabel metal3 s 177859 84328 178659 84448 6 i_dout0_1[7]
port 63 nsew signal input
rlabel metal2 s 148598 0 148654 800 6 i_dout0_1[8]
port 64 nsew signal input
rlabel metal3 s 177859 96160 178659 96280 6 i_dout0_1[9]
port 65 nsew signal input
rlabel metal2 s 570 180003 626 180803 6 io_in[0]
port 66 nsew signal input
rlabel metal2 s 36266 180003 36322 180803 6 io_in[10]
port 67 nsew signal input
rlabel metal2 s 39854 180003 39910 180803 6 io_in[11]
port 68 nsew signal input
rlabel metal2 s 43442 180003 43498 180803 6 io_in[12]
port 69 nsew signal input
rlabel metal2 s 46938 180003 46994 180803 6 io_in[13]
port 70 nsew signal input
rlabel metal2 s 50526 180003 50582 180803 6 io_in[14]
port 71 nsew signal input
rlabel metal2 s 54114 180003 54170 180803 6 io_in[15]
port 72 nsew signal input
rlabel metal2 s 57702 180003 57758 180803 6 io_in[16]
port 73 nsew signal input
rlabel metal2 s 61290 180003 61346 180803 6 io_in[17]
port 74 nsew signal input
rlabel metal2 s 64878 180003 64934 180803 6 io_in[18]
port 75 nsew signal input
rlabel metal2 s 68374 180003 68430 180803 6 io_in[19]
port 76 nsew signal input
rlabel metal2 s 4066 180003 4122 180803 6 io_in[1]
port 77 nsew signal input
rlabel metal2 s 71962 180003 72018 180803 6 io_in[20]
port 78 nsew signal input
rlabel metal2 s 75550 180003 75606 180803 6 io_in[21]
port 79 nsew signal input
rlabel metal2 s 79138 180003 79194 180803 6 io_in[22]
port 80 nsew signal input
rlabel metal2 s 82726 180003 82782 180803 6 io_in[23]
port 81 nsew signal input
rlabel metal2 s 86314 180003 86370 180803 6 io_in[24]
port 82 nsew signal input
rlabel metal2 s 89902 180003 89958 180803 6 io_in[25]
port 83 nsew signal input
rlabel metal2 s 93398 180003 93454 180803 6 io_in[26]
port 84 nsew signal input
rlabel metal2 s 96986 180003 97042 180803 6 io_in[27]
port 85 nsew signal input
rlabel metal2 s 100574 180003 100630 180803 6 io_in[28]
port 86 nsew signal input
rlabel metal2 s 104162 180003 104218 180803 6 io_in[29]
port 87 nsew signal input
rlabel metal2 s 7654 180003 7710 180803 6 io_in[2]
port 88 nsew signal input
rlabel metal2 s 107750 180003 107806 180803 6 io_in[30]
port 89 nsew signal input
rlabel metal2 s 111338 180003 111394 180803 6 io_in[31]
port 90 nsew signal input
rlabel metal2 s 114834 180003 114890 180803 6 io_in[32]
port 91 nsew signal input
rlabel metal2 s 118422 180003 118478 180803 6 io_in[33]
port 92 nsew signal input
rlabel metal2 s 122010 180003 122066 180803 6 io_in[34]
port 93 nsew signal input
rlabel metal2 s 125598 180003 125654 180803 6 io_in[35]
port 94 nsew signal input
rlabel metal2 s 129186 180003 129242 180803 6 io_in[36]
port 95 nsew signal input
rlabel metal2 s 132774 180003 132830 180803 6 io_in[37]
port 96 nsew signal input
rlabel metal2 s 11242 180003 11298 180803 6 io_in[3]
port 97 nsew signal input
rlabel metal2 s 14830 180003 14886 180803 6 io_in[4]
port 98 nsew signal input
rlabel metal2 s 18418 180003 18474 180803 6 io_in[5]
port 99 nsew signal input
rlabel metal2 s 22006 180003 22062 180803 6 io_in[6]
port 100 nsew signal input
rlabel metal2 s 25502 180003 25558 180803 6 io_in[7]
port 101 nsew signal input
rlabel metal2 s 29090 180003 29146 180803 6 io_in[8]
port 102 nsew signal input
rlabel metal2 s 32678 180003 32734 180803 6 io_in[9]
port 103 nsew signal input
rlabel metal2 s 1674 180003 1730 180803 6 io_oeb[0]
port 104 nsew signal output
rlabel metal2 s 37462 180003 37518 180803 6 io_oeb[10]
port 105 nsew signal output
rlabel metal2 s 41050 180003 41106 180803 6 io_oeb[11]
port 106 nsew signal output
rlabel metal2 s 44638 180003 44694 180803 6 io_oeb[12]
port 107 nsew signal output
rlabel metal2 s 48134 180003 48190 180803 6 io_oeb[13]
port 108 nsew signal output
rlabel metal2 s 51722 180003 51778 180803 6 io_oeb[14]
port 109 nsew signal output
rlabel metal2 s 55310 180003 55366 180803 6 io_oeb[15]
port 110 nsew signal output
rlabel metal2 s 58898 180003 58954 180803 6 io_oeb[16]
port 111 nsew signal output
rlabel metal2 s 62486 180003 62542 180803 6 io_oeb[17]
port 112 nsew signal output
rlabel metal2 s 66074 180003 66130 180803 6 io_oeb[18]
port 113 nsew signal output
rlabel metal2 s 69570 180003 69626 180803 6 io_oeb[19]
port 114 nsew signal output
rlabel metal2 s 5262 180003 5318 180803 6 io_oeb[1]
port 115 nsew signal output
rlabel metal2 s 73158 180003 73214 180803 6 io_oeb[20]
port 116 nsew signal output
rlabel metal2 s 76746 180003 76802 180803 6 io_oeb[21]
port 117 nsew signal output
rlabel metal2 s 80334 180003 80390 180803 6 io_oeb[22]
port 118 nsew signal output
rlabel metal2 s 83922 180003 83978 180803 6 io_oeb[23]
port 119 nsew signal output
rlabel metal2 s 87510 180003 87566 180803 6 io_oeb[24]
port 120 nsew signal output
rlabel metal2 s 91006 180003 91062 180803 6 io_oeb[25]
port 121 nsew signal output
rlabel metal2 s 94594 180003 94650 180803 6 io_oeb[26]
port 122 nsew signal output
rlabel metal2 s 98182 180003 98238 180803 6 io_oeb[27]
port 123 nsew signal output
rlabel metal2 s 101770 180003 101826 180803 6 io_oeb[28]
port 124 nsew signal output
rlabel metal2 s 105358 180003 105414 180803 6 io_oeb[29]
port 125 nsew signal output
rlabel metal2 s 8850 180003 8906 180803 6 io_oeb[2]
port 126 nsew signal output
rlabel metal2 s 108946 180003 109002 180803 6 io_oeb[30]
port 127 nsew signal output
rlabel metal2 s 112442 180003 112498 180803 6 io_oeb[31]
port 128 nsew signal output
rlabel metal2 s 116030 180003 116086 180803 6 io_oeb[32]
port 129 nsew signal output
rlabel metal2 s 119618 180003 119674 180803 6 io_oeb[33]
port 130 nsew signal output
rlabel metal2 s 123206 180003 123262 180803 6 io_oeb[34]
port 131 nsew signal output
rlabel metal2 s 126794 180003 126850 180803 6 io_oeb[35]
port 132 nsew signal output
rlabel metal2 s 130382 180003 130438 180803 6 io_oeb[36]
port 133 nsew signal output
rlabel metal2 s 133970 180003 134026 180803 6 io_oeb[37]
port 134 nsew signal output
rlabel metal2 s 12438 180003 12494 180803 6 io_oeb[3]
port 135 nsew signal output
rlabel metal2 s 16026 180003 16082 180803 6 io_oeb[4]
port 136 nsew signal output
rlabel metal2 s 19614 180003 19670 180803 6 io_oeb[5]
port 137 nsew signal output
rlabel metal2 s 23110 180003 23166 180803 6 io_oeb[6]
port 138 nsew signal output
rlabel metal2 s 26698 180003 26754 180803 6 io_oeb[7]
port 139 nsew signal output
rlabel metal2 s 30286 180003 30342 180803 6 io_oeb[8]
port 140 nsew signal output
rlabel metal2 s 33874 180003 33930 180803 6 io_oeb[9]
port 141 nsew signal output
rlabel metal2 s 2870 180003 2926 180803 6 io_out[0]
port 142 nsew signal output
rlabel metal2 s 38658 180003 38714 180803 6 io_out[10]
port 143 nsew signal output
rlabel metal2 s 42246 180003 42302 180803 6 io_out[11]
port 144 nsew signal output
rlabel metal2 s 45742 180003 45798 180803 6 io_out[12]
port 145 nsew signal output
rlabel metal2 s 49330 180003 49386 180803 6 io_out[13]
port 146 nsew signal output
rlabel metal2 s 52918 180003 52974 180803 6 io_out[14]
port 147 nsew signal output
rlabel metal2 s 56506 180003 56562 180803 6 io_out[15]
port 148 nsew signal output
rlabel metal2 s 60094 180003 60150 180803 6 io_out[16]
port 149 nsew signal output
rlabel metal2 s 63682 180003 63738 180803 6 io_out[17]
port 150 nsew signal output
rlabel metal2 s 67270 180003 67326 180803 6 io_out[18]
port 151 nsew signal output
rlabel metal2 s 70766 180003 70822 180803 6 io_out[19]
port 152 nsew signal output
rlabel metal2 s 6458 180003 6514 180803 6 io_out[1]
port 153 nsew signal output
rlabel metal2 s 74354 180003 74410 180803 6 io_out[20]
port 154 nsew signal output
rlabel metal2 s 77942 180003 77998 180803 6 io_out[21]
port 155 nsew signal output
rlabel metal2 s 81530 180003 81586 180803 6 io_out[22]
port 156 nsew signal output
rlabel metal2 s 85118 180003 85174 180803 6 io_out[23]
port 157 nsew signal output
rlabel metal2 s 88706 180003 88762 180803 6 io_out[24]
port 158 nsew signal output
rlabel metal2 s 92202 180003 92258 180803 6 io_out[25]
port 159 nsew signal output
rlabel metal2 s 95790 180003 95846 180803 6 io_out[26]
port 160 nsew signal output
rlabel metal2 s 99378 180003 99434 180803 6 io_out[27]
port 161 nsew signal output
rlabel metal2 s 102966 180003 103022 180803 6 io_out[28]
port 162 nsew signal output
rlabel metal2 s 106554 180003 106610 180803 6 io_out[29]
port 163 nsew signal output
rlabel metal2 s 10046 180003 10102 180803 6 io_out[2]
port 164 nsew signal output
rlabel metal2 s 110142 180003 110198 180803 6 io_out[30]
port 165 nsew signal output
rlabel metal2 s 113638 180003 113694 180803 6 io_out[31]
port 166 nsew signal output
rlabel metal2 s 117226 180003 117282 180803 6 io_out[32]
port 167 nsew signal output
rlabel metal2 s 120814 180003 120870 180803 6 io_out[33]
port 168 nsew signal output
rlabel metal2 s 124402 180003 124458 180803 6 io_out[34]
port 169 nsew signal output
rlabel metal2 s 127990 180003 128046 180803 6 io_out[35]
port 170 nsew signal output
rlabel metal2 s 131578 180003 131634 180803 6 io_out[36]
port 171 nsew signal output
rlabel metal2 s 135074 180003 135130 180803 6 io_out[37]
port 172 nsew signal output
rlabel metal2 s 13634 180003 13690 180803 6 io_out[3]
port 173 nsew signal output
rlabel metal2 s 17222 180003 17278 180803 6 io_out[4]
port 174 nsew signal output
rlabel metal2 s 20810 180003 20866 180803 6 io_out[5]
port 175 nsew signal output
rlabel metal2 s 24306 180003 24362 180803 6 io_out[6]
port 176 nsew signal output
rlabel metal2 s 27894 180003 27950 180803 6 io_out[7]
port 177 nsew signal output
rlabel metal2 s 31482 180003 31538 180803 6 io_out[8]
port 178 nsew signal output
rlabel metal2 s 35070 180003 35126 180803 6 io_out[9]
port 179 nsew signal output
rlabel metal2 s 130198 0 130254 800 6 irq[0]
port 180 nsew signal output
rlabel metal2 s 131486 0 131542 800 6 irq[1]
port 181 nsew signal output
rlabel metal2 s 132682 0 132738 800 6 irq[2]
port 182 nsew signal output
rlabel metal2 s 136270 180003 136326 180803 6 o_csb0
port 183 nsew signal output
rlabel metal2 s 135166 0 135222 800 6 o_csb0_1
port 184 nsew signal output
rlabel metal3 s 177859 9664 178659 9784 6 o_din0[0]
port 185 nsew signal output
rlabel metal2 s 154670 0 154726 800 6 o_din0[10]
port 186 nsew signal output
rlabel metal2 s 153014 180003 153070 180803 6 o_din0[11]
port 187 nsew signal output
rlabel metal3 s 0 85824 800 85944 6 o_din0[12]
port 188 nsew signal output
rlabel metal3 s 0 94664 800 94784 6 o_din0[13]
port 189 nsew signal output
rlabel metal2 s 159638 0 159694 800 6 o_din0[14]
port 190 nsew signal output
rlabel metal2 s 162030 0 162086 800 6 o_din0[15]
port 191 nsew signal output
rlabel metal3 s 177859 119688 178659 119808 6 o_din0[16]
port 192 nsew signal output
rlabel metal2 s 160098 180003 160154 180803 6 o_din0[17]
port 193 nsew signal output
rlabel metal3 s 0 107856 800 107976 6 o_din0[18]
port 194 nsew signal output
rlabel metal3 s 177859 135464 178659 135584 6 o_din0[19]
port 195 nsew signal output
rlabel metal2 s 137558 0 137614 800 6 o_din0[1]
port 196 nsew signal output
rlabel metal3 s 0 121184 800 121304 6 o_din0[20]
port 197 nsew signal output
rlabel metal3 s 0 130024 800 130144 6 o_din0[21]
port 198 nsew signal output
rlabel metal2 s 167274 180003 167330 180803 6 o_din0[22]
port 199 nsew signal output
rlabel metal3 s 177859 147160 178659 147280 6 o_din0[23]
port 200 nsew signal output
rlabel metal3 s 177859 155048 178659 155168 6 o_din0[24]
port 201 nsew signal output
rlabel metal3 s 0 147568 800 147688 6 o_din0[25]
port 202 nsew signal output
rlabel metal2 s 171874 0 171930 800 6 o_din0[26]
port 203 nsew signal output
rlabel metal3 s 177859 166880 178659 167000 6 o_din0[27]
port 204 nsew signal output
rlabel metal3 s 0 169600 800 169720 6 o_din0[28]
port 205 nsew signal output
rlabel metal3 s 177859 170824 178659 170944 6 o_din0[29]
port 206 nsew signal output
rlabel metal2 s 142250 180003 142306 180803 6 o_din0[2]
port 207 nsew signal output
rlabel metal3 s 177859 174768 178659 174888 6 o_din0[30]
port 208 nsew signal output
rlabel metal2 s 178038 180003 178094 180803 6 o_din0[31]
port 209 nsew signal output
rlabel metal3 s 177859 56856 178659 56976 6 o_din0[3]
port 210 nsew signal output
rlabel metal3 s 0 46248 800 46368 6 o_din0[4]
port 211 nsew signal output
rlabel metal3 s 177859 72632 178659 72752 6 o_din0[5]
port 212 nsew signal output
rlabel metal3 s 177859 80384 178659 80504 6 o_din0[6]
port 213 nsew signal output
rlabel metal3 s 0 63792 800 63912 6 o_din0[7]
port 214 nsew signal output
rlabel metal2 s 151082 0 151138 800 6 o_din0[8]
port 215 nsew signal output
rlabel metal3 s 0 77120 800 77240 6 o_din0[9]
port 216 nsew signal output
rlabel metal3 s 177859 13608 178659 13728 6 o_din0_1[0]
port 217 nsew signal output
rlabel metal2 s 153474 0 153530 800 6 o_din0_1[10]
port 218 nsew signal output
rlabel metal2 s 151818 180003 151874 180803 6 o_din0_1[11]
port 219 nsew signal output
rlabel metal2 s 157154 0 157210 800 6 o_din0_1[12]
port 220 nsew signal output
rlabel metal3 s 0 90312 800 90432 6 o_din0_1[13]
port 221 nsew signal output
rlabel metal2 s 157706 180003 157762 180803 6 o_din0_1[14]
port 222 nsew signal output
rlabel metal3 s 177859 115744 178659 115864 6 o_din0_1[15]
port 223 nsew signal output
rlabel metal2 s 164514 0 164570 800 6 o_din0_1[16]
port 224 nsew signal output
rlabel metal3 s 177859 123632 178659 123752 6 o_din0_1[17]
port 225 nsew signal output
rlabel metal3 s 0 103504 800 103624 6 o_din0_1[18]
port 226 nsew signal output
rlabel metal3 s 177859 131520 178659 131640 6 o_din0_1[19]
port 227 nsew signal output
rlabel metal2 s 138662 180003 138718 180803 6 o_din0_1[1]
port 228 nsew signal output
rlabel metal3 s 0 116696 800 116816 6 o_din0_1[20]
port 229 nsew signal output
rlabel metal2 s 166078 180003 166134 180803 6 o_din0_1[21]
port 230 nsew signal output
rlabel metal3 s 0 138728 800 138848 6 o_din0_1[22]
port 231 nsew signal output
rlabel metal3 s 177859 143352 178659 143472 6 o_din0_1[23]
port 232 nsew signal output
rlabel metal2 s 169666 180003 169722 180803 6 o_din0_1[24]
port 233 nsew signal output
rlabel metal2 s 170586 0 170642 800 6 o_din0_1[25]
port 234 nsew signal output
rlabel metal3 s 177859 162936 178659 163056 6 o_din0_1[26]
port 235 nsew signal output
rlabel metal2 s 175554 0 175610 800 6 o_din0_1[27]
port 236 nsew signal output
rlabel metal3 s 0 165248 800 165368 6 o_din0_1[28]
port 237 nsew signal output
rlabel metal2 s 176750 0 176806 800 6 o_din0_1[29]
port 238 nsew signal output
rlabel metal3 s 0 19728 800 19848 6 o_din0_1[2]
port 239 nsew signal output
rlabel metal2 s 175646 180003 175702 180803 6 o_din0_1[30]
port 240 nsew signal output
rlabel metal2 s 176842 180003 176898 180803 6 o_din0_1[31]
port 241 nsew signal output
rlabel metal3 s 177859 52912 178659 53032 6 o_din0_1[3]
port 242 nsew signal output
rlabel metal3 s 0 41760 800 41880 6 o_din0_1[4]
port 243 nsew signal output
rlabel metal2 s 143722 0 143778 800 6 o_din0_1[5]
port 244 nsew signal output
rlabel metal3 s 0 59440 800 59560 6 o_din0_1[6]
port 245 nsew signal output
rlabel metal3 s 177859 88272 178659 88392 6 o_din0_1[7]
port 246 nsew signal output
rlabel metal3 s 0 68280 800 68400 6 o_din0_1[8]
port 247 nsew signal output
rlabel metal2 s 150622 180003 150678 180803 6 o_din0_1[9]
port 248 nsew signal output
rlabel metal3 s 0 10888 800 11008 6 o_waddr0[0]
port 249 nsew signal output
rlabel metal3 s 177859 33328 178659 33448 6 o_waddr0[1]
port 250 nsew signal output
rlabel metal2 s 138846 0 138902 800 6 o_waddr0[2]
port 251 nsew signal output
rlabel metal3 s 0 32920 800 33040 6 o_waddr0[3]
port 252 nsew signal output
rlabel metal3 s 0 50600 800 50720 6 o_waddr0[4]
port 253 nsew signal output
rlabel metal2 s 144918 0 144974 800 6 o_waddr0[5]
port 254 nsew signal output
rlabel metal2 s 147402 0 147458 800 6 o_waddr0[6]
port 255 nsew signal output
rlabel metal2 s 148230 180003 148286 180803 6 o_waddr0[7]
port 256 nsew signal output
rlabel metal3 s 0 72632 800 72752 6 o_waddr0[8]
port 257 nsew signal output
rlabel metal2 s 136362 0 136418 800 6 o_waddr0_1[0]
port 258 nsew signal output
rlabel metal3 s 177859 29384 178659 29504 6 o_waddr0_1[1]
port 259 nsew signal output
rlabel metal2 s 143446 180003 143502 180803 6 o_waddr0_1[2]
port 260 nsew signal output
rlabel metal3 s 0 28568 800 28688 6 o_waddr0_1[3]
port 261 nsew signal output
rlabel metal3 s 177859 68688 178659 68808 6 o_waddr0_1[4]
port 262 nsew signal output
rlabel metal2 s 145838 180003 145894 180803 6 o_waddr0_1[5]
port 263 nsew signal output
rlabel metal2 s 146114 0 146170 800 6 o_waddr0_1[6]
port 264 nsew signal output
rlabel metal3 s 177859 92216 178659 92336 6 o_waddr0_1[7]
port 265 nsew signal output
rlabel metal2 s 149426 180003 149482 180803 6 o_waddr0_1[8]
port 266 nsew signal output
rlabel metal3 s 0 2184 800 2304 6 o_web0
port 267 nsew signal output
rlabel metal3 s 177859 1912 178659 2032 6 o_web0_1
port 268 nsew signal output
rlabel metal3 s 177859 17552 178659 17672 6 o_wmask0[0]
port 269 nsew signal output
rlabel metal2 s 141054 180003 141110 180803 6 o_wmask0[1]
port 270 nsew signal output
rlabel metal3 s 177859 45024 178659 45144 6 o_wmask0[2]
port 271 nsew signal output
rlabel metal3 s 0 37408 800 37528 6 o_wmask0[3]
port 272 nsew signal output
rlabel metal3 s 177859 21496 178659 21616 6 o_wmask0_1[0]
port 273 nsew signal output
rlabel metal2 s 139858 180003 139914 180803 6 o_wmask0_1[1]
port 274 nsew signal output
rlabel metal2 s 140042 0 140098 800 6 o_wmask0_1[2]
port 275 nsew signal output
rlabel metal3 s 177859 60800 178659 60920 6 o_wmask0_1[3]
port 276 nsew signal output
rlabel metal3 s 0 6536 800 6656 6 rst_i
port 277 nsew signal input
rlabel metal4 s 4208 2128 4528 178480 6 vccd1
port 278 nsew power input
rlabel metal4 s 34928 2128 35248 178480 6 vccd1
port 278 nsew power input
rlabel metal4 s 65648 2128 65968 178480 6 vccd1
port 278 nsew power input
rlabel metal4 s 96368 2128 96688 178480 6 vccd1
port 278 nsew power input
rlabel metal4 s 127088 2128 127408 178480 6 vccd1
port 278 nsew power input
rlabel metal4 s 157808 2128 158128 178480 6 vccd1
port 278 nsew power input
rlabel metal4 s 19568 2128 19888 178480 6 vssd1
port 279 nsew ground input
rlabel metal4 s 50288 2128 50608 178480 6 vssd1
port 279 nsew ground input
rlabel metal4 s 81008 2128 81328 178480 6 vssd1
port 279 nsew ground input
rlabel metal4 s 111728 2128 112048 178480 6 vssd1
port 279 nsew ground input
rlabel metal4 s 142448 2128 142768 178480 6 vssd1
port 279 nsew ground input
rlabel metal4 s 173168 2128 173488 178480 6 vssd1
port 279 nsew ground input
rlabel metal2 s 570 0 626 800 6 wb_clk_i
port 280 nsew signal input
rlabel metal2 s 1766 0 1822 800 6 wb_rst_i
port 281 nsew signal input
rlabel metal2 s 2962 0 3018 800 6 wbs_ack_o
port 282 nsew signal output
rlabel metal2 s 7838 0 7894 800 6 wbs_adr_i[0]
port 283 nsew signal input
rlabel metal2 s 49514 0 49570 800 6 wbs_adr_i[10]
port 284 nsew signal input
rlabel metal2 s 53102 0 53158 800 6 wbs_adr_i[11]
port 285 nsew signal input
rlabel metal2 s 56782 0 56838 800 6 wbs_adr_i[12]
port 286 nsew signal input
rlabel metal2 s 60462 0 60518 800 6 wbs_adr_i[13]
port 287 nsew signal input
rlabel metal2 s 64142 0 64198 800 6 wbs_adr_i[14]
port 288 nsew signal input
rlabel metal2 s 67822 0 67878 800 6 wbs_adr_i[15]
port 289 nsew signal input
rlabel metal2 s 71502 0 71558 800 6 wbs_adr_i[16]
port 290 nsew signal input
rlabel metal2 s 75182 0 75238 800 6 wbs_adr_i[17]
port 291 nsew signal input
rlabel metal2 s 78862 0 78918 800 6 wbs_adr_i[18]
port 292 nsew signal input
rlabel metal2 s 82542 0 82598 800 6 wbs_adr_i[19]
port 293 nsew signal input
rlabel metal2 s 12806 0 12862 800 6 wbs_adr_i[1]
port 294 nsew signal input
rlabel metal2 s 86222 0 86278 800 6 wbs_adr_i[20]
port 295 nsew signal input
rlabel metal2 s 89902 0 89958 800 6 wbs_adr_i[21]
port 296 nsew signal input
rlabel metal2 s 93490 0 93546 800 6 wbs_adr_i[22]
port 297 nsew signal input
rlabel metal2 s 97170 0 97226 800 6 wbs_adr_i[23]
port 298 nsew signal input
rlabel metal2 s 100850 0 100906 800 6 wbs_adr_i[24]
port 299 nsew signal input
rlabel metal2 s 104530 0 104586 800 6 wbs_adr_i[25]
port 300 nsew signal input
rlabel metal2 s 108210 0 108266 800 6 wbs_adr_i[26]
port 301 nsew signal input
rlabel metal2 s 111890 0 111946 800 6 wbs_adr_i[27]
port 302 nsew signal input
rlabel metal2 s 115570 0 115626 800 6 wbs_adr_i[28]
port 303 nsew signal input
rlabel metal2 s 119250 0 119306 800 6 wbs_adr_i[29]
port 304 nsew signal input
rlabel metal2 s 17682 0 17738 800 6 wbs_adr_i[2]
port 305 nsew signal input
rlabel metal2 s 122930 0 122986 800 6 wbs_adr_i[30]
port 306 nsew signal input
rlabel metal2 s 126610 0 126666 800 6 wbs_adr_i[31]
port 307 nsew signal input
rlabel metal2 s 22558 0 22614 800 6 wbs_adr_i[3]
port 308 nsew signal input
rlabel metal2 s 27434 0 27490 800 6 wbs_adr_i[4]
port 309 nsew signal input
rlabel metal2 s 31114 0 31170 800 6 wbs_adr_i[5]
port 310 nsew signal input
rlabel metal2 s 34794 0 34850 800 6 wbs_adr_i[6]
port 311 nsew signal input
rlabel metal2 s 38474 0 38530 800 6 wbs_adr_i[7]
port 312 nsew signal input
rlabel metal2 s 42154 0 42210 800 6 wbs_adr_i[8]
port 313 nsew signal input
rlabel metal2 s 45834 0 45890 800 6 wbs_adr_i[9]
port 314 nsew signal input
rlabel metal2 s 4158 0 4214 800 6 wbs_cyc_i
port 315 nsew signal input
rlabel metal2 s 9126 0 9182 800 6 wbs_dat_i[0]
port 316 nsew signal input
rlabel metal2 s 50710 0 50766 800 6 wbs_dat_i[10]
port 317 nsew signal input
rlabel metal2 s 54390 0 54446 800 6 wbs_dat_i[11]
port 318 nsew signal input
rlabel metal2 s 58070 0 58126 800 6 wbs_dat_i[12]
port 319 nsew signal input
rlabel metal2 s 61750 0 61806 800 6 wbs_dat_i[13]
port 320 nsew signal input
rlabel metal2 s 65338 0 65394 800 6 wbs_dat_i[14]
port 321 nsew signal input
rlabel metal2 s 69018 0 69074 800 6 wbs_dat_i[15]
port 322 nsew signal input
rlabel metal2 s 72698 0 72754 800 6 wbs_dat_i[16]
port 323 nsew signal input
rlabel metal2 s 76378 0 76434 800 6 wbs_dat_i[17]
port 324 nsew signal input
rlabel metal2 s 80058 0 80114 800 6 wbs_dat_i[18]
port 325 nsew signal input
rlabel metal2 s 83738 0 83794 800 6 wbs_dat_i[19]
port 326 nsew signal input
rlabel metal2 s 14002 0 14058 800 6 wbs_dat_i[1]
port 327 nsew signal input
rlabel metal2 s 87418 0 87474 800 6 wbs_dat_i[20]
port 328 nsew signal input
rlabel metal2 s 91098 0 91154 800 6 wbs_dat_i[21]
port 329 nsew signal input
rlabel metal2 s 94778 0 94834 800 6 wbs_dat_i[22]
port 330 nsew signal input
rlabel metal2 s 98458 0 98514 800 6 wbs_dat_i[23]
port 331 nsew signal input
rlabel metal2 s 102138 0 102194 800 6 wbs_dat_i[24]
port 332 nsew signal input
rlabel metal2 s 105726 0 105782 800 6 wbs_dat_i[25]
port 333 nsew signal input
rlabel metal2 s 109406 0 109462 800 6 wbs_dat_i[26]
port 334 nsew signal input
rlabel metal2 s 113086 0 113142 800 6 wbs_dat_i[27]
port 335 nsew signal input
rlabel metal2 s 116766 0 116822 800 6 wbs_dat_i[28]
port 336 nsew signal input
rlabel metal2 s 120446 0 120502 800 6 wbs_dat_i[29]
port 337 nsew signal input
rlabel metal2 s 18878 0 18934 800 6 wbs_dat_i[2]
port 338 nsew signal input
rlabel metal2 s 124126 0 124182 800 6 wbs_dat_i[30]
port 339 nsew signal input
rlabel metal2 s 127806 0 127862 800 6 wbs_dat_i[31]
port 340 nsew signal input
rlabel metal2 s 23754 0 23810 800 6 wbs_dat_i[3]
port 341 nsew signal input
rlabel metal2 s 28630 0 28686 800 6 wbs_dat_i[4]
port 342 nsew signal input
rlabel metal2 s 32310 0 32366 800 6 wbs_dat_i[5]
port 343 nsew signal input
rlabel metal2 s 35990 0 36046 800 6 wbs_dat_i[6]
port 344 nsew signal input
rlabel metal2 s 39670 0 39726 800 6 wbs_dat_i[7]
port 345 nsew signal input
rlabel metal2 s 43350 0 43406 800 6 wbs_dat_i[8]
port 346 nsew signal input
rlabel metal2 s 47030 0 47086 800 6 wbs_dat_i[9]
port 347 nsew signal input
rlabel metal2 s 10322 0 10378 800 6 wbs_dat_o[0]
port 348 nsew signal output
rlabel metal2 s 51906 0 51962 800 6 wbs_dat_o[10]
port 349 nsew signal output
rlabel metal2 s 55586 0 55642 800 6 wbs_dat_o[11]
port 350 nsew signal output
rlabel metal2 s 59266 0 59322 800 6 wbs_dat_o[12]
port 351 nsew signal output
rlabel metal2 s 62946 0 63002 800 6 wbs_dat_o[13]
port 352 nsew signal output
rlabel metal2 s 66626 0 66682 800 6 wbs_dat_o[14]
port 353 nsew signal output
rlabel metal2 s 70306 0 70362 800 6 wbs_dat_o[15]
port 354 nsew signal output
rlabel metal2 s 73986 0 74042 800 6 wbs_dat_o[16]
port 355 nsew signal output
rlabel metal2 s 77574 0 77630 800 6 wbs_dat_o[17]
port 356 nsew signal output
rlabel metal2 s 81254 0 81310 800 6 wbs_dat_o[18]
port 357 nsew signal output
rlabel metal2 s 84934 0 84990 800 6 wbs_dat_o[19]
port 358 nsew signal output
rlabel metal2 s 15198 0 15254 800 6 wbs_dat_o[1]
port 359 nsew signal output
rlabel metal2 s 88614 0 88670 800 6 wbs_dat_o[20]
port 360 nsew signal output
rlabel metal2 s 92294 0 92350 800 6 wbs_dat_o[21]
port 361 nsew signal output
rlabel metal2 s 95974 0 96030 800 6 wbs_dat_o[22]
port 362 nsew signal output
rlabel metal2 s 99654 0 99710 800 6 wbs_dat_o[23]
port 363 nsew signal output
rlabel metal2 s 103334 0 103390 800 6 wbs_dat_o[24]
port 364 nsew signal output
rlabel metal2 s 107014 0 107070 800 6 wbs_dat_o[25]
port 365 nsew signal output
rlabel metal2 s 110694 0 110750 800 6 wbs_dat_o[26]
port 366 nsew signal output
rlabel metal2 s 114374 0 114430 800 6 wbs_dat_o[27]
port 367 nsew signal output
rlabel metal2 s 117962 0 118018 800 6 wbs_dat_o[28]
port 368 nsew signal output
rlabel metal2 s 121642 0 121698 800 6 wbs_dat_o[29]
port 369 nsew signal output
rlabel metal2 s 20074 0 20130 800 6 wbs_dat_o[2]
port 370 nsew signal output
rlabel metal2 s 125322 0 125378 800 6 wbs_dat_o[30]
port 371 nsew signal output
rlabel metal2 s 129002 0 129058 800 6 wbs_dat_o[31]
port 372 nsew signal output
rlabel metal2 s 25042 0 25098 800 6 wbs_dat_o[3]
port 373 nsew signal output
rlabel metal2 s 29918 0 29974 800 6 wbs_dat_o[4]
port 374 nsew signal output
rlabel metal2 s 33598 0 33654 800 6 wbs_dat_o[5]
port 375 nsew signal output
rlabel metal2 s 37278 0 37334 800 6 wbs_dat_o[6]
port 376 nsew signal output
rlabel metal2 s 40866 0 40922 800 6 wbs_dat_o[7]
port 377 nsew signal output
rlabel metal2 s 44546 0 44602 800 6 wbs_dat_o[8]
port 378 nsew signal output
rlabel metal2 s 48226 0 48282 800 6 wbs_dat_o[9]
port 379 nsew signal output
rlabel metal2 s 11518 0 11574 800 6 wbs_sel_i[0]
port 380 nsew signal input
rlabel metal2 s 16394 0 16450 800 6 wbs_sel_i[1]
port 381 nsew signal input
rlabel metal2 s 21362 0 21418 800 6 wbs_sel_i[2]
port 382 nsew signal input
rlabel metal2 s 26238 0 26294 800 6 wbs_sel_i[3]
port 383 nsew signal input
rlabel metal2 s 5446 0 5502 800 6 wbs_stb_i
port 384 nsew signal input
rlabel metal2 s 6642 0 6698 800 6 wbs_we_i
port 385 nsew signal input
<< properties >>
string LEFclass BLOCK
string FIXED_BBOX 0 0 178659 180803
string LEFview TRUE
string GDS_FILE /project/openlane/user_proj/runs/user_proj/results/magic/user_proj.gds
string GDS_END 81548228
string GDS_START 1386298
<< end >>

