magic
tech sky130A
magscale 1 2
timestamp 1643956454
<< obsli1 >>
rect 1104 1717 197587 198033
<< obsm1 >>
rect 750 960 197599 198416
<< metal2 >>
rect 570 199469 626 200269
rect 1766 199469 1822 200269
rect 2962 199469 3018 200269
rect 4250 199469 4306 200269
rect 5446 199469 5502 200269
rect 6734 199469 6790 200269
rect 7930 199469 7986 200269
rect 9218 199469 9274 200269
rect 10414 199469 10470 200269
rect 11702 199469 11758 200269
rect 12898 199469 12954 200269
rect 14186 199469 14242 200269
rect 15382 199469 15438 200269
rect 16670 199469 16726 200269
rect 17866 199469 17922 200269
rect 19062 199469 19118 200269
rect 20350 199469 20406 200269
rect 21546 199469 21602 200269
rect 22834 199469 22890 200269
rect 24030 199469 24086 200269
rect 25318 199469 25374 200269
rect 26514 199469 26570 200269
rect 27802 199469 27858 200269
rect 28998 199469 29054 200269
rect 30286 199469 30342 200269
rect 31482 199469 31538 200269
rect 32770 199469 32826 200269
rect 33966 199469 34022 200269
rect 35162 199469 35218 200269
rect 36450 199469 36506 200269
rect 37646 199469 37702 200269
rect 38934 199469 38990 200269
rect 40130 199469 40186 200269
rect 41418 199469 41474 200269
rect 42614 199469 42670 200269
rect 43902 199469 43958 200269
rect 45098 199469 45154 200269
rect 46386 199469 46442 200269
rect 47582 199469 47638 200269
rect 48870 199469 48926 200269
rect 50066 199469 50122 200269
rect 51262 199469 51318 200269
rect 52550 199469 52606 200269
rect 53746 199469 53802 200269
rect 55034 199469 55090 200269
rect 56230 199469 56286 200269
rect 57518 199469 57574 200269
rect 58714 199469 58770 200269
rect 60002 199469 60058 200269
rect 61198 199469 61254 200269
rect 62486 199469 62542 200269
rect 63682 199469 63738 200269
rect 64970 199469 65026 200269
rect 66166 199469 66222 200269
rect 67362 199469 67418 200269
rect 68650 199469 68706 200269
rect 69846 199469 69902 200269
rect 71134 199469 71190 200269
rect 72330 199469 72386 200269
rect 73618 199469 73674 200269
rect 74814 199469 74870 200269
rect 76102 199469 76158 200269
rect 77298 199469 77354 200269
rect 78586 199469 78642 200269
rect 79782 199469 79838 200269
rect 81070 199469 81126 200269
rect 82266 199469 82322 200269
rect 83462 199469 83518 200269
rect 84750 199469 84806 200269
rect 85946 199469 86002 200269
rect 87234 199469 87290 200269
rect 88430 199469 88486 200269
rect 89718 199469 89774 200269
rect 90914 199469 90970 200269
rect 92202 199469 92258 200269
rect 93398 199469 93454 200269
rect 94686 199469 94742 200269
rect 95882 199469 95938 200269
rect 97170 199469 97226 200269
rect 98366 199469 98422 200269
rect 99654 199469 99710 200269
rect 100850 199469 100906 200269
rect 102046 199469 102102 200269
rect 103334 199469 103390 200269
rect 104530 199469 104586 200269
rect 105818 199469 105874 200269
rect 107014 199469 107070 200269
rect 108302 199469 108358 200269
rect 109498 199469 109554 200269
rect 110786 199469 110842 200269
rect 111982 199469 112038 200269
rect 113270 199469 113326 200269
rect 114466 199469 114522 200269
rect 115754 199469 115810 200269
rect 116950 199469 117006 200269
rect 118146 199469 118202 200269
rect 119434 199469 119490 200269
rect 120630 199469 120686 200269
rect 121918 199469 121974 200269
rect 123114 199469 123170 200269
rect 124402 199469 124458 200269
rect 125598 199469 125654 200269
rect 126886 199469 126942 200269
rect 128082 199469 128138 200269
rect 129370 199469 129426 200269
rect 130566 199469 130622 200269
rect 131854 199469 131910 200269
rect 133050 199469 133106 200269
rect 134246 199469 134302 200269
rect 135534 199469 135590 200269
rect 136730 199469 136786 200269
rect 138018 199469 138074 200269
rect 139214 199469 139270 200269
rect 140502 199469 140558 200269
rect 141698 199469 141754 200269
rect 142986 199469 143042 200269
rect 144182 199469 144238 200269
rect 145470 199469 145526 200269
rect 146666 199469 146722 200269
rect 147954 199469 148010 200269
rect 149150 199469 149206 200269
rect 150346 199469 150402 200269
rect 151634 199469 151690 200269
rect 152830 199469 152886 200269
rect 154118 199469 154174 200269
rect 155314 199469 155370 200269
rect 156602 199469 156658 200269
rect 157798 199469 157854 200269
rect 159086 199469 159142 200269
rect 160282 199469 160338 200269
rect 161570 199469 161626 200269
rect 162766 199469 162822 200269
rect 164054 199469 164110 200269
rect 165250 199469 165306 200269
rect 166446 199469 166502 200269
rect 167734 199469 167790 200269
rect 168930 199469 168986 200269
rect 170218 199469 170274 200269
rect 171414 199469 171470 200269
rect 172702 199469 172758 200269
rect 173898 199469 173954 200269
rect 175186 199469 175242 200269
rect 176382 199469 176438 200269
rect 177670 199469 177726 200269
rect 178866 199469 178922 200269
rect 180154 199469 180210 200269
rect 181350 199469 181406 200269
rect 182546 199469 182602 200269
rect 183834 199469 183890 200269
rect 185030 199469 185086 200269
rect 186318 199469 186374 200269
rect 187514 199469 187570 200269
rect 188802 199469 188858 200269
rect 189998 199469 190054 200269
rect 191286 199469 191342 200269
rect 192482 199469 192538 200269
rect 193770 199469 193826 200269
rect 194966 199469 195022 200269
rect 196254 199469 196310 200269
rect 197450 199469 197506 200269
rect 754 0 810 800
rect 2226 0 2282 800
rect 3698 0 3754 800
rect 5170 0 5226 800
rect 6642 0 6698 800
rect 8114 0 8170 800
rect 9586 0 9642 800
rect 11058 0 11114 800
rect 12530 0 12586 800
rect 14002 0 14058 800
rect 15474 0 15530 800
rect 16946 0 17002 800
rect 18418 0 18474 800
rect 19890 0 19946 800
rect 21454 0 21510 800
rect 22926 0 22982 800
rect 24398 0 24454 800
rect 25870 0 25926 800
rect 27342 0 27398 800
rect 28814 0 28870 800
rect 30286 0 30342 800
rect 31758 0 31814 800
rect 33230 0 33286 800
rect 34702 0 34758 800
rect 36174 0 36230 800
rect 37646 0 37702 800
rect 39118 0 39174 800
rect 40682 0 40738 800
rect 42154 0 42210 800
rect 43626 0 43682 800
rect 45098 0 45154 800
rect 46570 0 46626 800
rect 48042 0 48098 800
rect 49514 0 49570 800
rect 50986 0 51042 800
rect 52458 0 52514 800
rect 53930 0 53986 800
rect 55402 0 55458 800
rect 56874 0 56930 800
rect 58346 0 58402 800
rect 59818 0 59874 800
rect 61382 0 61438 800
rect 62854 0 62910 800
rect 64326 0 64382 800
rect 65798 0 65854 800
rect 67270 0 67326 800
rect 68742 0 68798 800
rect 70214 0 70270 800
rect 71686 0 71742 800
rect 73158 0 73214 800
rect 74630 0 74686 800
rect 76102 0 76158 800
rect 77574 0 77630 800
rect 79046 0 79102 800
rect 80610 0 80666 800
rect 82082 0 82138 800
rect 83554 0 83610 800
rect 85026 0 85082 800
rect 86498 0 86554 800
rect 87970 0 88026 800
rect 89442 0 89498 800
rect 90914 0 90970 800
rect 92386 0 92442 800
rect 93858 0 93914 800
rect 95330 0 95386 800
rect 96802 0 96858 800
rect 98274 0 98330 800
rect 99838 0 99894 800
rect 101310 0 101366 800
rect 102782 0 102838 800
rect 104254 0 104310 800
rect 105726 0 105782 800
rect 107198 0 107254 800
rect 108670 0 108726 800
rect 110142 0 110198 800
rect 111614 0 111670 800
rect 113086 0 113142 800
rect 114558 0 114614 800
rect 116030 0 116086 800
rect 117502 0 117558 800
rect 118974 0 119030 800
rect 120538 0 120594 800
rect 122010 0 122066 800
rect 123482 0 123538 800
rect 124954 0 125010 800
rect 126426 0 126482 800
rect 127898 0 127954 800
rect 129370 0 129426 800
rect 130842 0 130898 800
rect 132314 0 132370 800
rect 133786 0 133842 800
rect 135258 0 135314 800
rect 136730 0 136786 800
rect 138202 0 138258 800
rect 139766 0 139822 800
rect 141238 0 141294 800
rect 142710 0 142766 800
rect 144182 0 144238 800
rect 145654 0 145710 800
rect 147126 0 147182 800
rect 148598 0 148654 800
rect 150070 0 150126 800
rect 151542 0 151598 800
rect 153014 0 153070 800
rect 154486 0 154542 800
rect 155958 0 156014 800
rect 157430 0 157486 800
rect 158902 0 158958 800
rect 160466 0 160522 800
rect 161938 0 161994 800
rect 163410 0 163466 800
rect 164882 0 164938 800
rect 166354 0 166410 800
rect 167826 0 167882 800
rect 169298 0 169354 800
rect 170770 0 170826 800
rect 172242 0 172298 800
rect 173714 0 173770 800
rect 175186 0 175242 800
rect 176658 0 176714 800
rect 178130 0 178186 800
rect 179694 0 179750 800
rect 181166 0 181222 800
rect 182638 0 182694 800
rect 184110 0 184166 800
rect 185582 0 185638 800
rect 187054 0 187110 800
rect 188526 0 188582 800
rect 189998 0 190054 800
rect 191470 0 191526 800
rect 192942 0 192998 800
rect 194414 0 194470 800
rect 195886 0 195942 800
rect 197358 0 197414 800
<< obsm2 >>
rect 756 199413 1710 199469
rect 1878 199413 2906 199469
rect 3074 199413 4194 199469
rect 4362 199413 5390 199469
rect 5558 199413 6678 199469
rect 6846 199413 7874 199469
rect 8042 199413 9162 199469
rect 9330 199413 10358 199469
rect 10526 199413 11646 199469
rect 11814 199413 12842 199469
rect 13010 199413 14130 199469
rect 14298 199413 15326 199469
rect 15494 199413 16614 199469
rect 16782 199413 17810 199469
rect 17978 199413 19006 199469
rect 19174 199413 20294 199469
rect 20462 199413 21490 199469
rect 21658 199413 22778 199469
rect 22946 199413 23974 199469
rect 24142 199413 25262 199469
rect 25430 199413 26458 199469
rect 26626 199413 27746 199469
rect 27914 199413 28942 199469
rect 29110 199413 30230 199469
rect 30398 199413 31426 199469
rect 31594 199413 32714 199469
rect 32882 199413 33910 199469
rect 34078 199413 35106 199469
rect 35274 199413 36394 199469
rect 36562 199413 37590 199469
rect 37758 199413 38878 199469
rect 39046 199413 40074 199469
rect 40242 199413 41362 199469
rect 41530 199413 42558 199469
rect 42726 199413 43846 199469
rect 44014 199413 45042 199469
rect 45210 199413 46330 199469
rect 46498 199413 47526 199469
rect 47694 199413 48814 199469
rect 48982 199413 50010 199469
rect 50178 199413 51206 199469
rect 51374 199413 52494 199469
rect 52662 199413 53690 199469
rect 53858 199413 54978 199469
rect 55146 199413 56174 199469
rect 56342 199413 57462 199469
rect 57630 199413 58658 199469
rect 58826 199413 59946 199469
rect 60114 199413 61142 199469
rect 61310 199413 62430 199469
rect 62598 199413 63626 199469
rect 63794 199413 64914 199469
rect 65082 199413 66110 199469
rect 66278 199413 67306 199469
rect 67474 199413 68594 199469
rect 68762 199413 69790 199469
rect 69958 199413 71078 199469
rect 71246 199413 72274 199469
rect 72442 199413 73562 199469
rect 73730 199413 74758 199469
rect 74926 199413 76046 199469
rect 76214 199413 77242 199469
rect 77410 199413 78530 199469
rect 78698 199413 79726 199469
rect 79894 199413 81014 199469
rect 81182 199413 82210 199469
rect 82378 199413 83406 199469
rect 83574 199413 84694 199469
rect 84862 199413 85890 199469
rect 86058 199413 87178 199469
rect 87346 199413 88374 199469
rect 88542 199413 89662 199469
rect 89830 199413 90858 199469
rect 91026 199413 92146 199469
rect 92314 199413 93342 199469
rect 93510 199413 94630 199469
rect 94798 199413 95826 199469
rect 95994 199413 97114 199469
rect 97282 199413 98310 199469
rect 98478 199413 99598 199469
rect 99766 199413 100794 199469
rect 100962 199413 101990 199469
rect 102158 199413 103278 199469
rect 103446 199413 104474 199469
rect 104642 199413 105762 199469
rect 105930 199413 106958 199469
rect 107126 199413 108246 199469
rect 108414 199413 109442 199469
rect 109610 199413 110730 199469
rect 110898 199413 111926 199469
rect 112094 199413 113214 199469
rect 113382 199413 114410 199469
rect 114578 199413 115698 199469
rect 115866 199413 116894 199469
rect 117062 199413 118090 199469
rect 118258 199413 119378 199469
rect 119546 199413 120574 199469
rect 120742 199413 121862 199469
rect 122030 199413 123058 199469
rect 123226 199413 124346 199469
rect 124514 199413 125542 199469
rect 125710 199413 126830 199469
rect 126998 199413 128026 199469
rect 128194 199413 129314 199469
rect 129482 199413 130510 199469
rect 130678 199413 131798 199469
rect 131966 199413 132994 199469
rect 133162 199413 134190 199469
rect 134358 199413 135478 199469
rect 135646 199413 136674 199469
rect 136842 199413 137962 199469
rect 138130 199413 139158 199469
rect 139326 199413 140446 199469
rect 140614 199413 141642 199469
rect 141810 199413 142930 199469
rect 143098 199413 144126 199469
rect 144294 199413 145414 199469
rect 145582 199413 146610 199469
rect 146778 199413 147898 199469
rect 148066 199413 149094 199469
rect 149262 199413 150290 199469
rect 150458 199413 151578 199469
rect 151746 199413 152774 199469
rect 152942 199413 154062 199469
rect 154230 199413 155258 199469
rect 155426 199413 156546 199469
rect 156714 199413 157742 199469
rect 157910 199413 159030 199469
rect 159198 199413 160226 199469
rect 160394 199413 161514 199469
rect 161682 199413 162710 199469
rect 162878 199413 163998 199469
rect 164166 199413 165194 199469
rect 165362 199413 166390 199469
rect 166558 199413 167678 199469
rect 167846 199413 168874 199469
rect 169042 199413 170162 199469
rect 170330 199413 171358 199469
rect 171526 199413 172646 199469
rect 172814 199413 173842 199469
rect 174010 199413 175130 199469
rect 175298 199413 176326 199469
rect 176494 199413 177614 199469
rect 177782 199413 178810 199469
rect 178978 199413 180098 199469
rect 180266 199413 181294 199469
rect 181462 199413 182490 199469
rect 182658 199413 183778 199469
rect 183946 199413 184974 199469
rect 185142 199413 186262 199469
rect 186430 199413 187458 199469
rect 187626 199413 188746 199469
rect 188914 199413 189942 199469
rect 190110 199413 191230 199469
rect 191398 199413 192426 199469
rect 192594 199413 193714 199469
rect 193882 199413 194910 199469
rect 195078 199413 196198 199469
rect 196366 199413 197394 199469
rect 756 856 197506 199413
rect 866 734 2170 856
rect 2338 734 3642 856
rect 3810 734 5114 856
rect 5282 734 6586 856
rect 6754 734 8058 856
rect 8226 734 9530 856
rect 9698 734 11002 856
rect 11170 734 12474 856
rect 12642 734 13946 856
rect 14114 734 15418 856
rect 15586 734 16890 856
rect 17058 734 18362 856
rect 18530 734 19834 856
rect 20002 734 21398 856
rect 21566 734 22870 856
rect 23038 734 24342 856
rect 24510 734 25814 856
rect 25982 734 27286 856
rect 27454 734 28758 856
rect 28926 734 30230 856
rect 30398 734 31702 856
rect 31870 734 33174 856
rect 33342 734 34646 856
rect 34814 734 36118 856
rect 36286 734 37590 856
rect 37758 734 39062 856
rect 39230 734 40626 856
rect 40794 734 42098 856
rect 42266 734 43570 856
rect 43738 734 45042 856
rect 45210 734 46514 856
rect 46682 734 47986 856
rect 48154 734 49458 856
rect 49626 734 50930 856
rect 51098 734 52402 856
rect 52570 734 53874 856
rect 54042 734 55346 856
rect 55514 734 56818 856
rect 56986 734 58290 856
rect 58458 734 59762 856
rect 59930 734 61326 856
rect 61494 734 62798 856
rect 62966 734 64270 856
rect 64438 734 65742 856
rect 65910 734 67214 856
rect 67382 734 68686 856
rect 68854 734 70158 856
rect 70326 734 71630 856
rect 71798 734 73102 856
rect 73270 734 74574 856
rect 74742 734 76046 856
rect 76214 734 77518 856
rect 77686 734 78990 856
rect 79158 734 80554 856
rect 80722 734 82026 856
rect 82194 734 83498 856
rect 83666 734 84970 856
rect 85138 734 86442 856
rect 86610 734 87914 856
rect 88082 734 89386 856
rect 89554 734 90858 856
rect 91026 734 92330 856
rect 92498 734 93802 856
rect 93970 734 95274 856
rect 95442 734 96746 856
rect 96914 734 98218 856
rect 98386 734 99782 856
rect 99950 734 101254 856
rect 101422 734 102726 856
rect 102894 734 104198 856
rect 104366 734 105670 856
rect 105838 734 107142 856
rect 107310 734 108614 856
rect 108782 734 110086 856
rect 110254 734 111558 856
rect 111726 734 113030 856
rect 113198 734 114502 856
rect 114670 734 115974 856
rect 116142 734 117446 856
rect 117614 734 118918 856
rect 119086 734 120482 856
rect 120650 734 121954 856
rect 122122 734 123426 856
rect 123594 734 124898 856
rect 125066 734 126370 856
rect 126538 734 127842 856
rect 128010 734 129314 856
rect 129482 734 130786 856
rect 130954 734 132258 856
rect 132426 734 133730 856
rect 133898 734 135202 856
rect 135370 734 136674 856
rect 136842 734 138146 856
rect 138314 734 139710 856
rect 139878 734 141182 856
rect 141350 734 142654 856
rect 142822 734 144126 856
rect 144294 734 145598 856
rect 145766 734 147070 856
rect 147238 734 148542 856
rect 148710 734 150014 856
rect 150182 734 151486 856
rect 151654 734 152958 856
rect 153126 734 154430 856
rect 154598 734 155902 856
rect 156070 734 157374 856
rect 157542 734 158846 856
rect 159014 734 160410 856
rect 160578 734 161882 856
rect 162050 734 163354 856
rect 163522 734 164826 856
rect 164994 734 166298 856
rect 166466 734 167770 856
rect 167938 734 169242 856
rect 169410 734 170714 856
rect 170882 734 172186 856
rect 172354 734 173658 856
rect 173826 734 175130 856
rect 175298 734 176602 856
rect 176770 734 178074 856
rect 178242 734 179638 856
rect 179806 734 181110 856
rect 181278 734 182582 856
rect 182750 734 184054 856
rect 184222 734 185526 856
rect 185694 734 186998 856
rect 187166 734 188470 856
rect 188638 734 189942 856
rect 190110 734 191414 856
rect 191582 734 192886 856
rect 193054 734 194358 856
rect 194526 734 195830 856
rect 195998 734 197302 856
rect 197470 734 197506 856
<< metal3 >>
rect 0 198024 800 198144
rect 197325 197752 198125 197872
rect 0 193808 800 193928
rect 197325 192992 198125 193112
rect 0 189456 800 189576
rect 197325 188232 198125 188352
rect 0 185240 800 185360
rect 197325 183472 198125 183592
rect 0 181024 800 181144
rect 197325 178712 198125 178832
rect 0 176672 800 176792
rect 197325 173952 198125 174072
rect 0 172456 800 172576
rect 197325 169192 198125 169312
rect 0 168240 800 168360
rect 197325 164432 198125 164552
rect 0 163888 800 164008
rect 0 159672 800 159792
rect 197325 159672 198125 159792
rect 0 155456 800 155576
rect 197325 154912 198125 155032
rect 0 151104 800 151224
rect 197325 150152 198125 150272
rect 0 146888 800 147008
rect 197325 145392 198125 145512
rect 0 142672 800 142792
rect 197325 140632 198125 140752
rect 0 138320 800 138440
rect 197325 135872 198125 135992
rect 0 134104 800 134224
rect 197325 130976 198125 131096
rect 0 129888 800 130008
rect 197325 126216 198125 126336
rect 0 125536 800 125656
rect 0 121320 800 121440
rect 197325 121456 198125 121576
rect 0 117104 800 117224
rect 197325 116696 198125 116816
rect 0 112752 800 112872
rect 197325 111936 198125 112056
rect 0 108536 800 108656
rect 197325 107176 198125 107296
rect 0 104320 800 104440
rect 197325 102416 198125 102536
rect 0 99968 800 100088
rect 197325 97656 198125 97776
rect 0 95752 800 95872
rect 197325 92896 198125 93016
rect 0 91536 800 91656
rect 197325 88136 198125 88256
rect 0 87184 800 87304
rect 197325 83376 198125 83496
rect 0 82968 800 83088
rect 0 78752 800 78872
rect 197325 78616 198125 78736
rect 0 74400 800 74520
rect 197325 73856 198125 73976
rect 0 70184 800 70304
rect 197325 69096 198125 69216
rect 0 65968 800 66088
rect 197325 64200 198125 64320
rect 0 61616 800 61736
rect 197325 59440 198125 59560
rect 0 57400 800 57520
rect 197325 54680 198125 54800
rect 0 53184 800 53304
rect 197325 49920 198125 50040
rect 0 48832 800 48952
rect 197325 45160 198125 45280
rect 0 44616 800 44736
rect 0 40400 800 40520
rect 197325 40400 198125 40520
rect 0 36048 800 36168
rect 197325 35640 198125 35760
rect 0 31832 800 31952
rect 197325 30880 198125 31000
rect 0 27616 800 27736
rect 197325 26120 198125 26240
rect 0 23264 800 23384
rect 197325 21360 198125 21480
rect 0 19048 800 19168
rect 197325 16600 198125 16720
rect 0 14832 800 14952
rect 197325 11840 198125 11960
rect 0 10480 800 10600
rect 197325 7080 198125 7200
rect 0 6264 800 6384
rect 197325 2320 198125 2440
rect 0 2048 800 2168
<< obsm3 >>
rect 880 197952 197511 198117
rect 880 197944 197245 197952
rect 800 197672 197245 197944
rect 800 194008 197511 197672
rect 880 193728 197511 194008
rect 800 193192 197511 193728
rect 800 192912 197245 193192
rect 800 189656 197511 192912
rect 880 189376 197511 189656
rect 800 188432 197511 189376
rect 800 188152 197245 188432
rect 800 185440 197511 188152
rect 880 185160 197511 185440
rect 800 183672 197511 185160
rect 800 183392 197245 183672
rect 800 181224 197511 183392
rect 880 180944 197511 181224
rect 800 178912 197511 180944
rect 800 178632 197245 178912
rect 800 176872 197511 178632
rect 880 176592 197511 176872
rect 800 174152 197511 176592
rect 800 173872 197245 174152
rect 800 172656 197511 173872
rect 880 172376 197511 172656
rect 800 169392 197511 172376
rect 800 169112 197245 169392
rect 800 168440 197511 169112
rect 880 168160 197511 168440
rect 800 164632 197511 168160
rect 800 164352 197245 164632
rect 800 164088 197511 164352
rect 880 163808 197511 164088
rect 800 159872 197511 163808
rect 880 159592 197245 159872
rect 800 155656 197511 159592
rect 880 155376 197511 155656
rect 800 155112 197511 155376
rect 800 154832 197245 155112
rect 800 151304 197511 154832
rect 880 151024 197511 151304
rect 800 150352 197511 151024
rect 800 150072 197245 150352
rect 800 147088 197511 150072
rect 880 146808 197511 147088
rect 800 145592 197511 146808
rect 800 145312 197245 145592
rect 800 142872 197511 145312
rect 880 142592 197511 142872
rect 800 140832 197511 142592
rect 800 140552 197245 140832
rect 800 138520 197511 140552
rect 880 138240 197511 138520
rect 800 136072 197511 138240
rect 800 135792 197245 136072
rect 800 134304 197511 135792
rect 880 134024 197511 134304
rect 800 131176 197511 134024
rect 800 130896 197245 131176
rect 800 130088 197511 130896
rect 880 129808 197511 130088
rect 800 126416 197511 129808
rect 800 126136 197245 126416
rect 800 125736 197511 126136
rect 880 125456 197511 125736
rect 800 121656 197511 125456
rect 800 121520 197245 121656
rect 880 121376 197245 121520
rect 880 121240 197511 121376
rect 800 117304 197511 121240
rect 880 117024 197511 117304
rect 800 116896 197511 117024
rect 800 116616 197245 116896
rect 800 112952 197511 116616
rect 880 112672 197511 112952
rect 800 112136 197511 112672
rect 800 111856 197245 112136
rect 800 108736 197511 111856
rect 880 108456 197511 108736
rect 800 107376 197511 108456
rect 800 107096 197245 107376
rect 800 104520 197511 107096
rect 880 104240 197511 104520
rect 800 102616 197511 104240
rect 800 102336 197245 102616
rect 800 100168 197511 102336
rect 880 99888 197511 100168
rect 800 97856 197511 99888
rect 800 97576 197245 97856
rect 800 95952 197511 97576
rect 880 95672 197511 95952
rect 800 93096 197511 95672
rect 800 92816 197245 93096
rect 800 91736 197511 92816
rect 880 91456 197511 91736
rect 800 88336 197511 91456
rect 800 88056 197245 88336
rect 800 87384 197511 88056
rect 880 87104 197511 87384
rect 800 83576 197511 87104
rect 800 83296 197245 83576
rect 800 83168 197511 83296
rect 880 82888 197511 83168
rect 800 78952 197511 82888
rect 880 78816 197511 78952
rect 880 78672 197245 78816
rect 800 78536 197245 78672
rect 800 74600 197511 78536
rect 880 74320 197511 74600
rect 800 74056 197511 74320
rect 800 73776 197245 74056
rect 800 70384 197511 73776
rect 880 70104 197511 70384
rect 800 69296 197511 70104
rect 800 69016 197245 69296
rect 800 66168 197511 69016
rect 880 65888 197511 66168
rect 800 64400 197511 65888
rect 800 64120 197245 64400
rect 800 61816 197511 64120
rect 880 61536 197511 61816
rect 800 59640 197511 61536
rect 800 59360 197245 59640
rect 800 57600 197511 59360
rect 880 57320 197511 57600
rect 800 54880 197511 57320
rect 800 54600 197245 54880
rect 800 53384 197511 54600
rect 880 53104 197511 53384
rect 800 50120 197511 53104
rect 800 49840 197245 50120
rect 800 49032 197511 49840
rect 880 48752 197511 49032
rect 800 45360 197511 48752
rect 800 45080 197245 45360
rect 800 44816 197511 45080
rect 880 44536 197511 44816
rect 800 40600 197511 44536
rect 880 40320 197245 40600
rect 800 36248 197511 40320
rect 880 35968 197511 36248
rect 800 35840 197511 35968
rect 800 35560 197245 35840
rect 800 32032 197511 35560
rect 880 31752 197511 32032
rect 800 31080 197511 31752
rect 800 30800 197245 31080
rect 800 27816 197511 30800
rect 880 27536 197511 27816
rect 800 26320 197511 27536
rect 800 26040 197245 26320
rect 800 23464 197511 26040
rect 880 23184 197511 23464
rect 800 21560 197511 23184
rect 800 21280 197245 21560
rect 800 19248 197511 21280
rect 880 18968 197511 19248
rect 800 16800 197511 18968
rect 800 16520 197245 16800
rect 800 15032 197511 16520
rect 880 14752 197511 15032
rect 800 12040 197511 14752
rect 800 11760 197245 12040
rect 800 10680 197511 11760
rect 880 10400 197511 10680
rect 800 7280 197511 10400
rect 800 7000 197245 7280
rect 800 6464 197511 7000
rect 880 6184 197511 6464
rect 800 2520 197511 6184
rect 800 2248 197245 2520
rect 880 2240 197245 2248
rect 880 1968 197511 2240
rect 800 1803 197511 1968
<< metal4 >>
rect 4208 2128 4528 198064
rect 19568 2128 19888 198064
rect 34928 2128 35248 198064
rect 50288 2128 50608 198064
rect 65648 2128 65968 198064
rect 81008 2128 81328 198064
rect 96368 2128 96688 198064
rect 111728 2128 112048 198064
rect 127088 2128 127408 198064
rect 142448 2128 142768 198064
rect 157808 2128 158128 198064
rect 173168 2128 173488 198064
rect 188528 2128 188848 198064
<< obsm4 >>
rect 19195 3979 19488 197845
rect 19968 3979 34848 197845
rect 35328 3979 50208 197845
rect 50688 3979 65568 197845
rect 66048 3979 80928 197845
rect 81408 3979 96288 197845
rect 96768 3979 111648 197845
rect 112128 3979 127008 197845
rect 127488 3979 142368 197845
rect 142848 3979 157728 197845
rect 158208 3979 173088 197845
rect 173568 3979 188448 197845
rect 188928 3979 195901 197845
<< labels >>
rlabel metal2 s 141698 199469 141754 200269 6 clk_i
port 1 nsew signal input
rlabel metal2 s 145470 199469 145526 200269 6 i_dout0[0]
port 2 nsew signal input
rlabel metal3 s 0 82968 800 83088 6 i_dout0[10]
port 3 nsew signal input
rlabel metal3 s 0 91536 800 91656 6 i_dout0[11]
port 4 nsew signal input
rlabel metal2 s 166446 199469 166502 200269 6 i_dout0[12]
port 5 nsew signal input
rlabel metal3 s 0 104320 800 104440 6 i_dout0[13]
port 6 nsew signal input
rlabel metal2 s 181166 0 181222 800 6 i_dout0[14]
port 7 nsew signal input
rlabel metal2 s 182638 0 182694 800 6 i_dout0[15]
port 8 nsew signal input
rlabel metal3 s 0 117104 800 117224 6 i_dout0[16]
port 9 nsew signal input
rlabel metal2 s 172702 199469 172758 200269 6 i_dout0[17]
port 10 nsew signal input
rlabel metal2 s 175186 199469 175242 200269 6 i_dout0[18]
port 11 nsew signal input
rlabel metal3 s 197325 159672 198125 159792 6 i_dout0[19]
port 12 nsew signal input
rlabel metal3 s 0 14832 800 14952 6 i_dout0[1]
port 13 nsew signal input
rlabel metal3 s 0 138320 800 138440 6 i_dout0[20]
port 14 nsew signal input
rlabel metal2 s 185582 0 185638 800 6 i_dout0[21]
port 15 nsew signal input
rlabel metal3 s 197325 164432 198125 164552 6 i_dout0[22]
port 16 nsew signal input
rlabel metal3 s 0 155456 800 155576 6 i_dout0[23]
port 17 nsew signal input
rlabel metal2 s 189998 0 190054 800 6 i_dout0[24]
port 18 nsew signal input
rlabel metal2 s 186318 199469 186374 200269 6 i_dout0[25]
port 19 nsew signal input
rlabel metal3 s 0 176672 800 176792 6 i_dout0[26]
port 20 nsew signal input
rlabel metal3 s 0 181024 800 181144 6 i_dout0[27]
port 21 nsew signal input
rlabel metal3 s 197325 183472 198125 183592 6 i_dout0[28]
port 22 nsew signal input
rlabel metal2 s 195886 0 195942 800 6 i_dout0[29]
port 23 nsew signal input
rlabel metal3 s 197325 35640 198125 35760 6 i_dout0[2]
port 24 nsew signal input
rlabel metal2 s 194966 199469 195022 200269 6 i_dout0[30]
port 25 nsew signal input
rlabel metal2 s 197358 0 197414 800 6 i_dout0[31]
port 26 nsew signal input
rlabel metal3 s 0 40400 800 40520 6 i_dout0[3]
port 27 nsew signal input
rlabel metal3 s 0 48832 800 48952 6 i_dout0[4]
port 28 nsew signal input
rlabel metal2 s 173714 0 173770 800 6 i_dout0[5]
port 29 nsew signal input
rlabel metal3 s 197325 73856 198125 73976 6 i_dout0[6]
port 30 nsew signal input
rlabel metal3 s 197325 97656 198125 97776 6 i_dout0[7]
port 31 nsew signal input
rlabel metal2 s 160282 199469 160338 200269 6 i_dout0[8]
port 32 nsew signal input
rlabel metal3 s 0 74400 800 74520 6 i_dout0[9]
port 33 nsew signal input
rlabel metal2 s 163410 0 163466 800 6 i_dout0_1[0]
port 34 nsew signal input
rlabel metal3 s 197325 126216 198125 126336 6 i_dout0_1[10]
port 35 nsew signal input
rlabel metal3 s 0 87184 800 87304 6 i_dout0_1[11]
port 36 nsew signal input
rlabel metal2 s 165250 199469 165306 200269 6 i_dout0_1[12]
port 37 nsew signal input
rlabel metal2 s 178130 0 178186 800 6 i_dout0_1[13]
port 38 nsew signal input
rlabel metal3 s 197325 135872 198125 135992 6 i_dout0_1[14]
port 39 nsew signal input
rlabel metal2 s 168930 199469 168986 200269 6 i_dout0_1[15]
port 40 nsew signal input
rlabel metal2 s 171414 199469 171470 200269 6 i_dout0_1[16]
port 41 nsew signal input
rlabel metal3 s 0 121320 800 121440 6 i_dout0_1[17]
port 42 nsew signal input
rlabel metal2 s 173898 199469 173954 200269 6 i_dout0_1[18]
port 43 nsew signal input
rlabel metal2 s 176382 199469 176438 200269 6 i_dout0_1[19]
port 44 nsew signal input
rlabel metal2 s 164882 0 164938 800 6 i_dout0_1[1]
port 45 nsew signal input
rlabel metal3 s 0 134104 800 134224 6 i_dout0_1[20]
port 46 nsew signal input
rlabel metal2 s 181350 199469 181406 200269 6 i_dout0_1[21]
port 47 nsew signal input
rlabel metal2 s 187054 0 187110 800 6 i_dout0_1[22]
port 48 nsew signal input
rlabel metal3 s 0 151104 800 151224 6 i_dout0_1[23]
port 49 nsew signal input
rlabel metal2 s 185030 199469 185086 200269 6 i_dout0_1[24]
port 50 nsew signal input
rlabel metal3 s 197325 173952 198125 174072 6 i_dout0_1[25]
port 51 nsew signal input
rlabel metal2 s 191470 0 191526 800 6 i_dout0_1[26]
port 52 nsew signal input
rlabel metal3 s 197325 178712 198125 178832 6 i_dout0_1[27]
port 53 nsew signal input
rlabel metal2 s 191286 199469 191342 200269 6 i_dout0_1[28]
port 54 nsew signal input
rlabel metal3 s 197325 188232 198125 188352 6 i_dout0_1[29]
port 55 nsew signal input
rlabel metal3 s 197325 30880 198125 31000 6 i_dout0_1[2]
port 56 nsew signal input
rlabel metal2 s 193770 199469 193826 200269 6 i_dout0_1[30]
port 57 nsew signal input
rlabel metal3 s 0 193808 800 193928 6 i_dout0_1[31]
port 58 nsew signal input
rlabel metal3 s 197325 45160 198125 45280 6 i_dout0_1[3]
port 59 nsew signal input
rlabel metal3 s 0 44616 800 44736 6 i_dout0_1[4]
port 60 nsew signal input
rlabel metal2 s 152830 199469 152886 200269 6 i_dout0_1[5]
port 61 nsew signal input
rlabel metal2 s 155314 199469 155370 200269 6 i_dout0_1[6]
port 62 nsew signal input
rlabel metal3 s 197325 92896 198125 93016 6 i_dout0_1[7]
port 63 nsew signal input
rlabel metal2 s 159086 199469 159142 200269 6 i_dout0_1[8]
port 64 nsew signal input
rlabel metal3 s 197325 121456 198125 121576 6 i_dout0_1[9]
port 65 nsew signal input
rlabel metal2 s 570 199469 626 200269 6 io_in[0]
port 66 nsew signal input
rlabel metal2 s 37646 199469 37702 200269 6 io_in[10]
port 67 nsew signal input
rlabel metal2 s 41418 199469 41474 200269 6 io_in[11]
port 68 nsew signal input
rlabel metal2 s 45098 199469 45154 200269 6 io_in[12]
port 69 nsew signal input
rlabel metal2 s 48870 199469 48926 200269 6 io_in[13]
port 70 nsew signal input
rlabel metal2 s 52550 199469 52606 200269 6 io_in[14]
port 71 nsew signal input
rlabel metal2 s 56230 199469 56286 200269 6 io_in[15]
port 72 nsew signal input
rlabel metal2 s 60002 199469 60058 200269 6 io_in[16]
port 73 nsew signal input
rlabel metal2 s 63682 199469 63738 200269 6 io_in[17]
port 74 nsew signal input
rlabel metal2 s 67362 199469 67418 200269 6 io_in[18]
port 75 nsew signal input
rlabel metal2 s 71134 199469 71190 200269 6 io_in[19]
port 76 nsew signal input
rlabel metal2 s 4250 199469 4306 200269 6 io_in[1]
port 77 nsew signal input
rlabel metal2 s 74814 199469 74870 200269 6 io_in[20]
port 78 nsew signal input
rlabel metal2 s 78586 199469 78642 200269 6 io_in[21]
port 79 nsew signal input
rlabel metal2 s 82266 199469 82322 200269 6 io_in[22]
port 80 nsew signal input
rlabel metal2 s 85946 199469 86002 200269 6 io_in[23]
port 81 nsew signal input
rlabel metal2 s 89718 199469 89774 200269 6 io_in[24]
port 82 nsew signal input
rlabel metal2 s 93398 199469 93454 200269 6 io_in[25]
port 83 nsew signal input
rlabel metal2 s 97170 199469 97226 200269 6 io_in[26]
port 84 nsew signal input
rlabel metal2 s 100850 199469 100906 200269 6 io_in[27]
port 85 nsew signal input
rlabel metal2 s 104530 199469 104586 200269 6 io_in[28]
port 86 nsew signal input
rlabel metal2 s 108302 199469 108358 200269 6 io_in[29]
port 87 nsew signal input
rlabel metal2 s 7930 199469 7986 200269 6 io_in[2]
port 88 nsew signal input
rlabel metal2 s 111982 199469 112038 200269 6 io_in[30]
port 89 nsew signal input
rlabel metal2 s 115754 199469 115810 200269 6 io_in[31]
port 90 nsew signal input
rlabel metal2 s 119434 199469 119490 200269 6 io_in[32]
port 91 nsew signal input
rlabel metal2 s 123114 199469 123170 200269 6 io_in[33]
port 92 nsew signal input
rlabel metal2 s 126886 199469 126942 200269 6 io_in[34]
port 93 nsew signal input
rlabel metal2 s 130566 199469 130622 200269 6 io_in[35]
port 94 nsew signal input
rlabel metal2 s 134246 199469 134302 200269 6 io_in[36]
port 95 nsew signal input
rlabel metal2 s 138018 199469 138074 200269 6 io_in[37]
port 96 nsew signal input
rlabel metal2 s 11702 199469 11758 200269 6 io_in[3]
port 97 nsew signal input
rlabel metal2 s 15382 199469 15438 200269 6 io_in[4]
port 98 nsew signal input
rlabel metal2 s 19062 199469 19118 200269 6 io_in[5]
port 99 nsew signal input
rlabel metal2 s 22834 199469 22890 200269 6 io_in[6]
port 100 nsew signal input
rlabel metal2 s 26514 199469 26570 200269 6 io_in[7]
port 101 nsew signal input
rlabel metal2 s 30286 199469 30342 200269 6 io_in[8]
port 102 nsew signal input
rlabel metal2 s 33966 199469 34022 200269 6 io_in[9]
port 103 nsew signal input
rlabel metal2 s 1766 199469 1822 200269 6 io_oeb[0]
port 104 nsew signal output
rlabel metal2 s 38934 199469 38990 200269 6 io_oeb[10]
port 105 nsew signal output
rlabel metal2 s 42614 199469 42670 200269 6 io_oeb[11]
port 106 nsew signal output
rlabel metal2 s 46386 199469 46442 200269 6 io_oeb[12]
port 107 nsew signal output
rlabel metal2 s 50066 199469 50122 200269 6 io_oeb[13]
port 108 nsew signal output
rlabel metal2 s 53746 199469 53802 200269 6 io_oeb[14]
port 109 nsew signal output
rlabel metal2 s 57518 199469 57574 200269 6 io_oeb[15]
port 110 nsew signal output
rlabel metal2 s 61198 199469 61254 200269 6 io_oeb[16]
port 111 nsew signal output
rlabel metal2 s 64970 199469 65026 200269 6 io_oeb[17]
port 112 nsew signal output
rlabel metal2 s 68650 199469 68706 200269 6 io_oeb[18]
port 113 nsew signal output
rlabel metal2 s 72330 199469 72386 200269 6 io_oeb[19]
port 114 nsew signal output
rlabel metal2 s 5446 199469 5502 200269 6 io_oeb[1]
port 115 nsew signal output
rlabel metal2 s 76102 199469 76158 200269 6 io_oeb[20]
port 116 nsew signal output
rlabel metal2 s 79782 199469 79838 200269 6 io_oeb[21]
port 117 nsew signal output
rlabel metal2 s 83462 199469 83518 200269 6 io_oeb[22]
port 118 nsew signal output
rlabel metal2 s 87234 199469 87290 200269 6 io_oeb[23]
port 119 nsew signal output
rlabel metal2 s 90914 199469 90970 200269 6 io_oeb[24]
port 120 nsew signal output
rlabel metal2 s 94686 199469 94742 200269 6 io_oeb[25]
port 121 nsew signal output
rlabel metal2 s 98366 199469 98422 200269 6 io_oeb[26]
port 122 nsew signal output
rlabel metal2 s 102046 199469 102102 200269 6 io_oeb[27]
port 123 nsew signal output
rlabel metal2 s 105818 199469 105874 200269 6 io_oeb[28]
port 124 nsew signal output
rlabel metal2 s 109498 199469 109554 200269 6 io_oeb[29]
port 125 nsew signal output
rlabel metal2 s 9218 199469 9274 200269 6 io_oeb[2]
port 126 nsew signal output
rlabel metal2 s 113270 199469 113326 200269 6 io_oeb[30]
port 127 nsew signal output
rlabel metal2 s 116950 199469 117006 200269 6 io_oeb[31]
port 128 nsew signal output
rlabel metal2 s 120630 199469 120686 200269 6 io_oeb[32]
port 129 nsew signal output
rlabel metal2 s 124402 199469 124458 200269 6 io_oeb[33]
port 130 nsew signal output
rlabel metal2 s 128082 199469 128138 200269 6 io_oeb[34]
port 131 nsew signal output
rlabel metal2 s 131854 199469 131910 200269 6 io_oeb[35]
port 132 nsew signal output
rlabel metal2 s 135534 199469 135590 200269 6 io_oeb[36]
port 133 nsew signal output
rlabel metal2 s 139214 199469 139270 200269 6 io_oeb[37]
port 134 nsew signal output
rlabel metal2 s 12898 199469 12954 200269 6 io_oeb[3]
port 135 nsew signal output
rlabel metal2 s 16670 199469 16726 200269 6 io_oeb[4]
port 136 nsew signal output
rlabel metal2 s 20350 199469 20406 200269 6 io_oeb[5]
port 137 nsew signal output
rlabel metal2 s 24030 199469 24086 200269 6 io_oeb[6]
port 138 nsew signal output
rlabel metal2 s 27802 199469 27858 200269 6 io_oeb[7]
port 139 nsew signal output
rlabel metal2 s 31482 199469 31538 200269 6 io_oeb[8]
port 140 nsew signal output
rlabel metal2 s 35162 199469 35218 200269 6 io_oeb[9]
port 141 nsew signal output
rlabel metal2 s 2962 199469 3018 200269 6 io_out[0]
port 142 nsew signal output
rlabel metal2 s 40130 199469 40186 200269 6 io_out[10]
port 143 nsew signal output
rlabel metal2 s 43902 199469 43958 200269 6 io_out[11]
port 144 nsew signal output
rlabel metal2 s 47582 199469 47638 200269 6 io_out[12]
port 145 nsew signal output
rlabel metal2 s 51262 199469 51318 200269 6 io_out[13]
port 146 nsew signal output
rlabel metal2 s 55034 199469 55090 200269 6 io_out[14]
port 147 nsew signal output
rlabel metal2 s 58714 199469 58770 200269 6 io_out[15]
port 148 nsew signal output
rlabel metal2 s 62486 199469 62542 200269 6 io_out[16]
port 149 nsew signal output
rlabel metal2 s 66166 199469 66222 200269 6 io_out[17]
port 150 nsew signal output
rlabel metal2 s 69846 199469 69902 200269 6 io_out[18]
port 151 nsew signal output
rlabel metal2 s 73618 199469 73674 200269 6 io_out[19]
port 152 nsew signal output
rlabel metal2 s 6734 199469 6790 200269 6 io_out[1]
port 153 nsew signal output
rlabel metal2 s 77298 199469 77354 200269 6 io_out[20]
port 154 nsew signal output
rlabel metal2 s 81070 199469 81126 200269 6 io_out[21]
port 155 nsew signal output
rlabel metal2 s 84750 199469 84806 200269 6 io_out[22]
port 156 nsew signal output
rlabel metal2 s 88430 199469 88486 200269 6 io_out[23]
port 157 nsew signal output
rlabel metal2 s 92202 199469 92258 200269 6 io_out[24]
port 158 nsew signal output
rlabel metal2 s 95882 199469 95938 200269 6 io_out[25]
port 159 nsew signal output
rlabel metal2 s 99654 199469 99710 200269 6 io_out[26]
port 160 nsew signal output
rlabel metal2 s 103334 199469 103390 200269 6 io_out[27]
port 161 nsew signal output
rlabel metal2 s 107014 199469 107070 200269 6 io_out[28]
port 162 nsew signal output
rlabel metal2 s 110786 199469 110842 200269 6 io_out[29]
port 163 nsew signal output
rlabel metal2 s 10414 199469 10470 200269 6 io_out[2]
port 164 nsew signal output
rlabel metal2 s 114466 199469 114522 200269 6 io_out[30]
port 165 nsew signal output
rlabel metal2 s 118146 199469 118202 200269 6 io_out[31]
port 166 nsew signal output
rlabel metal2 s 121918 199469 121974 200269 6 io_out[32]
port 167 nsew signal output
rlabel metal2 s 125598 199469 125654 200269 6 io_out[33]
port 168 nsew signal output
rlabel metal2 s 129370 199469 129426 200269 6 io_out[34]
port 169 nsew signal output
rlabel metal2 s 133050 199469 133106 200269 6 io_out[35]
port 170 nsew signal output
rlabel metal2 s 136730 199469 136786 200269 6 io_out[36]
port 171 nsew signal output
rlabel metal2 s 140502 199469 140558 200269 6 io_out[37]
port 172 nsew signal output
rlabel metal2 s 14186 199469 14242 200269 6 io_out[3]
port 173 nsew signal output
rlabel metal2 s 17866 199469 17922 200269 6 io_out[4]
port 174 nsew signal output
rlabel metal2 s 21546 199469 21602 200269 6 io_out[5]
port 175 nsew signal output
rlabel metal2 s 25318 199469 25374 200269 6 io_out[6]
port 176 nsew signal output
rlabel metal2 s 28998 199469 29054 200269 6 io_out[7]
port 177 nsew signal output
rlabel metal2 s 32770 199469 32826 200269 6 io_out[8]
port 178 nsew signal output
rlabel metal2 s 36450 199469 36506 200269 6 io_out[9]
port 179 nsew signal output
rlabel metal2 s 157430 0 157486 800 6 irq[0]
port 180 nsew signal output
rlabel metal2 s 158902 0 158958 800 6 irq[1]
port 181 nsew signal output
rlabel metal2 s 160466 0 160522 800 6 irq[2]
port 182 nsew signal output
rlabel metal2 s 142986 199469 143042 200269 6 o_csb0
port 183 nsew signal output
rlabel metal3 s 197325 2320 198125 2440 6 o_csb0_1
port 184 nsew signal output
rlabel metal2 s 146666 199469 146722 200269 6 o_din0[0]
port 185 nsew signal output
rlabel metal2 s 164054 199469 164110 200269 6 o_din0[10]
port 186 nsew signal output
rlabel metal3 s 0 95752 800 95872 6 o_din0[11]
port 187 nsew signal output
rlabel metal3 s 0 99968 800 100088 6 o_din0[12]
port 188 nsew signal output
rlabel metal2 s 179694 0 179750 800 6 o_din0[13]
port 189 nsew signal output
rlabel metal2 s 167734 199469 167790 200269 6 o_din0[14]
port 190 nsew signal output
rlabel metal3 s 197325 140632 198125 140752 6 o_din0[15]
port 191 nsew signal output
rlabel metal3 s 197325 150152 198125 150272 6 o_din0[16]
port 192 nsew signal output
rlabel metal3 s 0 125536 800 125656 6 o_din0[17]
port 193 nsew signal output
rlabel metal2 s 184110 0 184166 800 6 o_din0[18]
port 194 nsew signal output
rlabel metal2 s 178866 199469 178922 200269 6 o_din0[19]
port 195 nsew signal output
rlabel metal2 s 166354 0 166410 800 6 o_din0[1]
port 196 nsew signal output
rlabel metal2 s 180154 199469 180210 200269 6 o_din0[20]
port 197 nsew signal output
rlabel metal2 s 183834 199469 183890 200269 6 o_din0[21]
port 198 nsew signal output
rlabel metal3 s 0 146888 800 147008 6 o_din0[22]
port 199 nsew signal output
rlabel metal3 s 0 159672 800 159792 6 o_din0[23]
port 200 nsew signal output
rlabel metal3 s 0 168240 800 168360 6 o_din0[24]
port 201 nsew signal output
rlabel metal2 s 187514 199469 187570 200269 6 o_din0[25]
port 202 nsew signal output
rlabel metal2 s 192942 0 192998 800 6 o_din0[26]
port 203 nsew signal output
rlabel metal2 s 189998 199469 190054 200269 6 o_din0[27]
port 204 nsew signal output
rlabel metal2 s 194414 0 194470 800 6 o_din0[28]
port 205 nsew signal output
rlabel metal2 s 192482 199469 192538 200269 6 o_din0[29]
port 206 nsew signal output
rlabel metal3 s 0 31832 800 31952 6 o_din0[2]
port 207 nsew signal output
rlabel metal3 s 197325 197752 198125 197872 6 o_din0[30]
port 208 nsew signal output
rlabel metal2 s 197450 199469 197506 200269 6 o_din0[31]
port 209 nsew signal output
rlabel metal3 s 197325 49920 198125 50040 6 o_din0[3]
port 210 nsew signal output
rlabel metal3 s 0 57400 800 57520 6 o_din0[4]
port 211 nsew signal output
rlabel metal3 s 197325 69096 198125 69216 6 o_din0[5]
port 212 nsew signal output
rlabel metal2 s 156602 199469 156658 200269 6 o_din0[6]
port 213 nsew signal output
rlabel metal3 s 0 65968 800 66088 6 o_din0[7]
port 214 nsew signal output
rlabel metal3 s 197325 111936 198125 112056 6 o_din0[8]
port 215 nsew signal output
rlabel metal3 s 0 78752 800 78872 6 o_din0[9]
port 216 nsew signal output
rlabel metal3 s 0 6264 800 6384 6 o_din0_1[0]
port 217 nsew signal output
rlabel metal2 s 175186 0 175242 800 6 o_din0_1[10]
port 218 nsew signal output
rlabel metal3 s 197325 130976 198125 131096 6 o_din0_1[11]
port 219 nsew signal output
rlabel metal2 s 176658 0 176714 800 6 o_din0_1[12]
port 220 nsew signal output
rlabel metal3 s 0 108536 800 108656 6 o_din0_1[13]
port 221 nsew signal output
rlabel metal3 s 0 112752 800 112872 6 o_din0_1[14]
port 222 nsew signal output
rlabel metal2 s 170218 199469 170274 200269 6 o_din0_1[15]
port 223 nsew signal output
rlabel metal3 s 197325 145392 198125 145512 6 o_din0_1[16]
port 224 nsew signal output
rlabel metal3 s 197325 154912 198125 155032 6 o_din0_1[17]
port 225 nsew signal output
rlabel metal3 s 0 129888 800 130008 6 o_din0_1[18]
port 226 nsew signal output
rlabel metal2 s 177670 199469 177726 200269 6 o_din0_1[19]
port 227 nsew signal output
rlabel metal3 s 197325 21360 198125 21480 6 o_din0_1[1]
port 228 nsew signal output
rlabel metal3 s 0 142672 800 142792 6 o_din0_1[20]
port 229 nsew signal output
rlabel metal2 s 182546 199469 182602 200269 6 o_din0_1[21]
port 230 nsew signal output
rlabel metal2 s 188526 0 188582 800 6 o_din0_1[22]
port 231 nsew signal output
rlabel metal3 s 197325 169192 198125 169312 6 o_din0_1[23]
port 232 nsew signal output
rlabel metal3 s 0 163888 800 164008 6 o_din0_1[24]
port 233 nsew signal output
rlabel metal3 s 0 172456 800 172576 6 o_din0_1[25]
port 234 nsew signal output
rlabel metal2 s 188802 199469 188858 200269 6 o_din0_1[26]
port 235 nsew signal output
rlabel metal3 s 0 185240 800 185360 6 o_din0_1[27]
port 236 nsew signal output
rlabel metal3 s 0 189456 800 189576 6 o_din0_1[28]
port 237 nsew signal output
rlabel metal3 s 197325 192992 198125 193112 6 o_din0_1[29]
port 238 nsew signal output
rlabel metal2 s 147954 199469 148010 200269 6 o_din0_1[2]
port 239 nsew signal output
rlabel metal2 s 196254 199469 196310 200269 6 o_din0_1[30]
port 240 nsew signal output
rlabel metal3 s 0 198024 800 198144 6 o_din0_1[31]
port 241 nsew signal output
rlabel metal2 s 149150 199469 149206 200269 6 o_din0_1[3]
port 242 nsew signal output
rlabel metal3 s 0 53184 800 53304 6 o_din0_1[4]
port 243 nsew signal output
rlabel metal3 s 197325 64200 198125 64320 6 o_din0_1[5]
port 244 nsew signal output
rlabel metal3 s 197325 78616 198125 78736 6 o_din0_1[6]
port 245 nsew signal output
rlabel metal2 s 157798 199469 157854 200269 6 o_din0_1[7]
port 246 nsew signal output
rlabel metal3 s 197325 107176 198125 107296 6 o_din0_1[8]
port 247 nsew signal output
rlabel metal2 s 162766 199469 162822 200269 6 o_din0_1[9]
port 248 nsew signal output
rlabel metal3 s 197325 7080 198125 7200 6 o_waddr0[0]
port 249 nsew signal output
rlabel metal3 s 197325 26120 198125 26240 6 o_waddr0[1]
port 250 nsew signal output
rlabel metal2 s 167826 0 167882 800 6 o_waddr0[2]
port 251 nsew signal output
rlabel metal2 s 150346 199469 150402 200269 6 o_waddr0[3]
port 252 nsew signal output
rlabel metal2 s 151634 199469 151690 200269 6 o_waddr0[4]
port 253 nsew signal output
rlabel metal3 s 0 61616 800 61736 6 o_waddr0[5]
port 254 nsew signal output
rlabel metal3 s 197325 88136 198125 88256 6 o_waddr0[6]
port 255 nsew signal output
rlabel metal3 s 0 70184 800 70304 6 o_waddr0[7]
port 256 nsew signal output
rlabel metal3 s 197325 116696 198125 116816 6 o_waddr0[8]
port 257 nsew signal output
rlabel metal3 s 0 10480 800 10600 6 o_waddr0_1[0]
port 258 nsew signal output
rlabel metal3 s 0 19048 800 19168 6 o_waddr0_1[1]
port 259 nsew signal output
rlabel metal3 s 0 36048 800 36168 6 o_waddr0_1[2]
port 260 nsew signal output
rlabel metal2 s 170770 0 170826 800 6 o_waddr0_1[3]
port 261 nsew signal output
rlabel metal3 s 197325 59440 198125 59560 6 o_waddr0_1[4]
port 262 nsew signal output
rlabel metal2 s 154118 199469 154174 200269 6 o_waddr0_1[5]
port 263 nsew signal output
rlabel metal3 s 197325 83376 198125 83496 6 o_waddr0_1[6]
port 264 nsew signal output
rlabel metal3 s 197325 102416 198125 102536 6 o_waddr0_1[7]
port 265 nsew signal output
rlabel metal2 s 161570 199469 161626 200269 6 o_waddr0_1[8]
port 266 nsew signal output
rlabel metal3 s 0 2048 800 2168 6 o_web0
port 267 nsew signal output
rlabel metal2 s 144182 199469 144238 200269 6 o_web0_1
port 268 nsew signal output
rlabel metal3 s 197325 11840 198125 11960 6 o_wmask0[0]
port 269 nsew signal output
rlabel metal3 s 0 27616 800 27736 6 o_wmask0[1]
port 270 nsew signal output
rlabel metal2 s 169298 0 169354 800 6 o_wmask0[2]
port 271 nsew signal output
rlabel metal2 s 172242 0 172298 800 6 o_wmask0[3]
port 272 nsew signal output
rlabel metal3 s 197325 16600 198125 16720 6 o_wmask0_1[0]
port 273 nsew signal output
rlabel metal3 s 0 23264 800 23384 6 o_wmask0_1[1]
port 274 nsew signal output
rlabel metal3 s 197325 40400 198125 40520 6 o_wmask0_1[2]
port 275 nsew signal output
rlabel metal3 s 197325 54680 198125 54800 6 o_wmask0_1[3]
port 276 nsew signal output
rlabel metal2 s 161938 0 161994 800 6 rst_i
port 277 nsew signal input
rlabel metal4 s 4208 2128 4528 198064 6 vccd1
port 278 nsew power input
rlabel metal4 s 34928 2128 35248 198064 6 vccd1
port 278 nsew power input
rlabel metal4 s 65648 2128 65968 198064 6 vccd1
port 278 nsew power input
rlabel metal4 s 96368 2128 96688 198064 6 vccd1
port 278 nsew power input
rlabel metal4 s 127088 2128 127408 198064 6 vccd1
port 278 nsew power input
rlabel metal4 s 157808 2128 158128 198064 6 vccd1
port 278 nsew power input
rlabel metal4 s 188528 2128 188848 198064 6 vccd1
port 278 nsew power input
rlabel metal4 s 19568 2128 19888 198064 6 vssd1
port 279 nsew ground input
rlabel metal4 s 50288 2128 50608 198064 6 vssd1
port 279 nsew ground input
rlabel metal4 s 81008 2128 81328 198064 6 vssd1
port 279 nsew ground input
rlabel metal4 s 111728 2128 112048 198064 6 vssd1
port 279 nsew ground input
rlabel metal4 s 142448 2128 142768 198064 6 vssd1
port 279 nsew ground input
rlabel metal4 s 173168 2128 173488 198064 6 vssd1
port 279 nsew ground input
rlabel metal2 s 754 0 810 800 6 wb_clk_i
port 280 nsew signal input
rlabel metal2 s 2226 0 2282 800 6 wb_rst_i
port 281 nsew signal input
rlabel metal2 s 3698 0 3754 800 6 wbs_ack_o
port 282 nsew signal output
rlabel metal2 s 9586 0 9642 800 6 wbs_adr_i[0]
port 283 nsew signal input
rlabel metal2 s 59818 0 59874 800 6 wbs_adr_i[10]
port 284 nsew signal input
rlabel metal2 s 64326 0 64382 800 6 wbs_adr_i[11]
port 285 nsew signal input
rlabel metal2 s 68742 0 68798 800 6 wbs_adr_i[12]
port 286 nsew signal input
rlabel metal2 s 73158 0 73214 800 6 wbs_adr_i[13]
port 287 nsew signal input
rlabel metal2 s 77574 0 77630 800 6 wbs_adr_i[14]
port 288 nsew signal input
rlabel metal2 s 82082 0 82138 800 6 wbs_adr_i[15]
port 289 nsew signal input
rlabel metal2 s 86498 0 86554 800 6 wbs_adr_i[16]
port 290 nsew signal input
rlabel metal2 s 90914 0 90970 800 6 wbs_adr_i[17]
port 291 nsew signal input
rlabel metal2 s 95330 0 95386 800 6 wbs_adr_i[18]
port 292 nsew signal input
rlabel metal2 s 99838 0 99894 800 6 wbs_adr_i[19]
port 293 nsew signal input
rlabel metal2 s 15474 0 15530 800 6 wbs_adr_i[1]
port 294 nsew signal input
rlabel metal2 s 104254 0 104310 800 6 wbs_adr_i[20]
port 295 nsew signal input
rlabel metal2 s 108670 0 108726 800 6 wbs_adr_i[21]
port 296 nsew signal input
rlabel metal2 s 113086 0 113142 800 6 wbs_adr_i[22]
port 297 nsew signal input
rlabel metal2 s 117502 0 117558 800 6 wbs_adr_i[23]
port 298 nsew signal input
rlabel metal2 s 122010 0 122066 800 6 wbs_adr_i[24]
port 299 nsew signal input
rlabel metal2 s 126426 0 126482 800 6 wbs_adr_i[25]
port 300 nsew signal input
rlabel metal2 s 130842 0 130898 800 6 wbs_adr_i[26]
port 301 nsew signal input
rlabel metal2 s 135258 0 135314 800 6 wbs_adr_i[27]
port 302 nsew signal input
rlabel metal2 s 139766 0 139822 800 6 wbs_adr_i[28]
port 303 nsew signal input
rlabel metal2 s 144182 0 144238 800 6 wbs_adr_i[29]
port 304 nsew signal input
rlabel metal2 s 21454 0 21510 800 6 wbs_adr_i[2]
port 305 nsew signal input
rlabel metal2 s 148598 0 148654 800 6 wbs_adr_i[30]
port 306 nsew signal input
rlabel metal2 s 153014 0 153070 800 6 wbs_adr_i[31]
port 307 nsew signal input
rlabel metal2 s 27342 0 27398 800 6 wbs_adr_i[3]
port 308 nsew signal input
rlabel metal2 s 33230 0 33286 800 6 wbs_adr_i[4]
port 309 nsew signal input
rlabel metal2 s 37646 0 37702 800 6 wbs_adr_i[5]
port 310 nsew signal input
rlabel metal2 s 42154 0 42210 800 6 wbs_adr_i[6]
port 311 nsew signal input
rlabel metal2 s 46570 0 46626 800 6 wbs_adr_i[7]
port 312 nsew signal input
rlabel metal2 s 50986 0 51042 800 6 wbs_adr_i[8]
port 313 nsew signal input
rlabel metal2 s 55402 0 55458 800 6 wbs_adr_i[9]
port 314 nsew signal input
rlabel metal2 s 5170 0 5226 800 6 wbs_cyc_i
port 315 nsew signal input
rlabel metal2 s 11058 0 11114 800 6 wbs_dat_i[0]
port 316 nsew signal input
rlabel metal2 s 61382 0 61438 800 6 wbs_dat_i[10]
port 317 nsew signal input
rlabel metal2 s 65798 0 65854 800 6 wbs_dat_i[11]
port 318 nsew signal input
rlabel metal2 s 70214 0 70270 800 6 wbs_dat_i[12]
port 319 nsew signal input
rlabel metal2 s 74630 0 74686 800 6 wbs_dat_i[13]
port 320 nsew signal input
rlabel metal2 s 79046 0 79102 800 6 wbs_dat_i[14]
port 321 nsew signal input
rlabel metal2 s 83554 0 83610 800 6 wbs_dat_i[15]
port 322 nsew signal input
rlabel metal2 s 87970 0 88026 800 6 wbs_dat_i[16]
port 323 nsew signal input
rlabel metal2 s 92386 0 92442 800 6 wbs_dat_i[17]
port 324 nsew signal input
rlabel metal2 s 96802 0 96858 800 6 wbs_dat_i[18]
port 325 nsew signal input
rlabel metal2 s 101310 0 101366 800 6 wbs_dat_i[19]
port 326 nsew signal input
rlabel metal2 s 16946 0 17002 800 6 wbs_dat_i[1]
port 327 nsew signal input
rlabel metal2 s 105726 0 105782 800 6 wbs_dat_i[20]
port 328 nsew signal input
rlabel metal2 s 110142 0 110198 800 6 wbs_dat_i[21]
port 329 nsew signal input
rlabel metal2 s 114558 0 114614 800 6 wbs_dat_i[22]
port 330 nsew signal input
rlabel metal2 s 118974 0 119030 800 6 wbs_dat_i[23]
port 331 nsew signal input
rlabel metal2 s 123482 0 123538 800 6 wbs_dat_i[24]
port 332 nsew signal input
rlabel metal2 s 127898 0 127954 800 6 wbs_dat_i[25]
port 333 nsew signal input
rlabel metal2 s 132314 0 132370 800 6 wbs_dat_i[26]
port 334 nsew signal input
rlabel metal2 s 136730 0 136786 800 6 wbs_dat_i[27]
port 335 nsew signal input
rlabel metal2 s 141238 0 141294 800 6 wbs_dat_i[28]
port 336 nsew signal input
rlabel metal2 s 145654 0 145710 800 6 wbs_dat_i[29]
port 337 nsew signal input
rlabel metal2 s 22926 0 22982 800 6 wbs_dat_i[2]
port 338 nsew signal input
rlabel metal2 s 150070 0 150126 800 6 wbs_dat_i[30]
port 339 nsew signal input
rlabel metal2 s 154486 0 154542 800 6 wbs_dat_i[31]
port 340 nsew signal input
rlabel metal2 s 28814 0 28870 800 6 wbs_dat_i[3]
port 341 nsew signal input
rlabel metal2 s 34702 0 34758 800 6 wbs_dat_i[4]
port 342 nsew signal input
rlabel metal2 s 39118 0 39174 800 6 wbs_dat_i[5]
port 343 nsew signal input
rlabel metal2 s 43626 0 43682 800 6 wbs_dat_i[6]
port 344 nsew signal input
rlabel metal2 s 48042 0 48098 800 6 wbs_dat_i[7]
port 345 nsew signal input
rlabel metal2 s 52458 0 52514 800 6 wbs_dat_i[8]
port 346 nsew signal input
rlabel metal2 s 56874 0 56930 800 6 wbs_dat_i[9]
port 347 nsew signal input
rlabel metal2 s 12530 0 12586 800 6 wbs_dat_o[0]
port 348 nsew signal output
rlabel metal2 s 62854 0 62910 800 6 wbs_dat_o[10]
port 349 nsew signal output
rlabel metal2 s 67270 0 67326 800 6 wbs_dat_o[11]
port 350 nsew signal output
rlabel metal2 s 71686 0 71742 800 6 wbs_dat_o[12]
port 351 nsew signal output
rlabel metal2 s 76102 0 76158 800 6 wbs_dat_o[13]
port 352 nsew signal output
rlabel metal2 s 80610 0 80666 800 6 wbs_dat_o[14]
port 353 nsew signal output
rlabel metal2 s 85026 0 85082 800 6 wbs_dat_o[15]
port 354 nsew signal output
rlabel metal2 s 89442 0 89498 800 6 wbs_dat_o[16]
port 355 nsew signal output
rlabel metal2 s 93858 0 93914 800 6 wbs_dat_o[17]
port 356 nsew signal output
rlabel metal2 s 98274 0 98330 800 6 wbs_dat_o[18]
port 357 nsew signal output
rlabel metal2 s 102782 0 102838 800 6 wbs_dat_o[19]
port 358 nsew signal output
rlabel metal2 s 18418 0 18474 800 6 wbs_dat_o[1]
port 359 nsew signal output
rlabel metal2 s 107198 0 107254 800 6 wbs_dat_o[20]
port 360 nsew signal output
rlabel metal2 s 111614 0 111670 800 6 wbs_dat_o[21]
port 361 nsew signal output
rlabel metal2 s 116030 0 116086 800 6 wbs_dat_o[22]
port 362 nsew signal output
rlabel metal2 s 120538 0 120594 800 6 wbs_dat_o[23]
port 363 nsew signal output
rlabel metal2 s 124954 0 125010 800 6 wbs_dat_o[24]
port 364 nsew signal output
rlabel metal2 s 129370 0 129426 800 6 wbs_dat_o[25]
port 365 nsew signal output
rlabel metal2 s 133786 0 133842 800 6 wbs_dat_o[26]
port 366 nsew signal output
rlabel metal2 s 138202 0 138258 800 6 wbs_dat_o[27]
port 367 nsew signal output
rlabel metal2 s 142710 0 142766 800 6 wbs_dat_o[28]
port 368 nsew signal output
rlabel metal2 s 147126 0 147182 800 6 wbs_dat_o[29]
port 369 nsew signal output
rlabel metal2 s 24398 0 24454 800 6 wbs_dat_o[2]
port 370 nsew signal output
rlabel metal2 s 151542 0 151598 800 6 wbs_dat_o[30]
port 371 nsew signal output
rlabel metal2 s 155958 0 156014 800 6 wbs_dat_o[31]
port 372 nsew signal output
rlabel metal2 s 30286 0 30342 800 6 wbs_dat_o[3]
port 373 nsew signal output
rlabel metal2 s 36174 0 36230 800 6 wbs_dat_o[4]
port 374 nsew signal output
rlabel metal2 s 40682 0 40738 800 6 wbs_dat_o[5]
port 375 nsew signal output
rlabel metal2 s 45098 0 45154 800 6 wbs_dat_o[6]
port 376 nsew signal output
rlabel metal2 s 49514 0 49570 800 6 wbs_dat_o[7]
port 377 nsew signal output
rlabel metal2 s 53930 0 53986 800 6 wbs_dat_o[8]
port 378 nsew signal output
rlabel metal2 s 58346 0 58402 800 6 wbs_dat_o[9]
port 379 nsew signal output
rlabel metal2 s 14002 0 14058 800 6 wbs_sel_i[0]
port 380 nsew signal input
rlabel metal2 s 19890 0 19946 800 6 wbs_sel_i[1]
port 381 nsew signal input
rlabel metal2 s 25870 0 25926 800 6 wbs_sel_i[2]
port 382 nsew signal input
rlabel metal2 s 31758 0 31814 800 6 wbs_sel_i[3]
port 383 nsew signal input
rlabel metal2 s 6642 0 6698 800 6 wbs_stb_i
port 384 nsew signal input
rlabel metal2 s 8114 0 8170 800 6 wbs_we_i
port 385 nsew signal input
<< properties >>
string LEFclass BLOCK
string FIXED_BBOX 0 0 198125 200269
string LEFview TRUE
string GDS_FILE /home/roman/projects/opencircuitdesign/shuttle5/caravel_mpw/openlane/user_proj/runs/user_proj/results/magic/user_proj.gds
string GDS_END 96742068
string GDS_START 1460676
<< end >>

