magic
tech sky130A
magscale 1 2
timestamp 1645590684
<< locali >>
rect 202153 243899 202187 244137
rect 218989 243491 219023 243865
rect 219081 243355 219115 243797
rect 42199 241145 42349 241179
rect 43361 240159 43395 241077
rect 45937 240363 45971 241145
rect 49617 240431 49651 241145
rect 50905 240227 50939 241145
rect 53481 240499 53515 241145
rect 54585 240295 54619 241145
rect 54677 240839 54711 241145
rect 57161 240567 57195 241213
rect 83013 240771 83047 241077
rect 115949 240771 115983 241145
rect 180901 240635 180935 240873
rect 182097 240703 182131 240873
rect 50353 3859 50387 4029
rect 50261 3791 50295 3825
rect 50445 3791 50479 4029
rect 50261 3757 50479 3791
rect 69673 3315 69707 3757
rect 122297 3179 122331 3689
<< viali >>
rect 202153 244137 202187 244171
rect 202153 243865 202187 243899
rect 218989 243865 219023 243899
rect 218989 243457 219023 243491
rect 219081 243797 219115 243831
rect 219081 243321 219115 243355
rect 57161 241213 57195 241247
rect 42165 241145 42199 241179
rect 42349 241145 42383 241179
rect 45937 241145 45971 241179
rect 43361 241077 43395 241111
rect 49617 241145 49651 241179
rect 49617 240397 49651 240431
rect 50905 241145 50939 241179
rect 45937 240329 45971 240363
rect 53481 241145 53515 241179
rect 53481 240465 53515 240499
rect 54585 241145 54619 241179
rect 54677 241145 54711 241179
rect 54677 240805 54711 240839
rect 115949 241145 115983 241179
rect 83013 241077 83047 241111
rect 83013 240737 83047 240771
rect 115949 240737 115983 240771
rect 180901 240873 180935 240907
rect 182097 240873 182131 240907
rect 182097 240669 182131 240703
rect 180901 240601 180935 240635
rect 57161 240533 57195 240567
rect 54585 240261 54619 240295
rect 50905 240193 50939 240227
rect 43361 240125 43395 240159
rect 50353 4029 50387 4063
rect 50261 3825 50295 3859
rect 50353 3825 50387 3859
rect 50445 4029 50479 4063
rect 69673 3757 69707 3791
rect 69673 3281 69707 3315
rect 122297 3689 122331 3723
rect 122297 3145 122331 3179
<< metal1 >>
rect 201494 702992 201500 703044
rect 201552 703032 201558 703044
rect 202782 703032 202788 703044
rect 201552 703004 202788 703032
rect 201552 702992 201558 703004
rect 202782 702992 202788 703004
rect 202840 702992 202846 703044
rect 333238 700612 333244 700664
rect 333296 700652 333302 700664
rect 364978 700652 364984 700664
rect 333296 700624 364984 700652
rect 333296 700612 333302 700624
rect 364978 700612 364984 700624
rect 365036 700612 365042 700664
rect 327718 700544 327724 700596
rect 327776 700584 327782 700596
rect 429838 700584 429844 700596
rect 327776 700556 429844 700584
rect 327776 700544 327782 700556
rect 429838 700544 429844 700556
rect 429896 700544 429902 700596
rect 330478 700476 330484 700528
rect 330536 700516 330542 700528
rect 462314 700516 462320 700528
rect 330536 700488 462320 700516
rect 330536 700476 330542 700488
rect 462314 700476 462320 700488
rect 462372 700476 462378 700528
rect 211798 700408 211804 700460
rect 211856 700448 211862 700460
rect 348786 700448 348792 700460
rect 211856 700420 348792 700448
rect 211856 700408 211862 700420
rect 348786 700408 348792 700420
rect 348844 700408 348850 700460
rect 105446 700340 105452 700392
rect 105504 700380 105510 700392
rect 106182 700380 106188 700392
rect 105504 700352 106188 700380
rect 105504 700340 105510 700352
rect 106182 700340 106188 700352
rect 106240 700340 106246 700392
rect 170306 700340 170312 700392
rect 170364 700380 170370 700392
rect 178034 700380 178040 700392
rect 170364 700352 178040 700380
rect 170364 700340 170370 700352
rect 178034 700340 178040 700352
rect 178092 700340 178098 700392
rect 193858 700340 193864 700392
rect 193916 700380 193922 700392
rect 332502 700380 332508 700392
rect 193916 700352 332508 700380
rect 193916 700340 193922 700352
rect 332502 700340 332508 700352
rect 332560 700340 332566 700392
rect 334618 700340 334624 700392
rect 334676 700380 334682 700392
rect 397454 700380 397460 700392
rect 334676 700352 397460 700380
rect 334676 700340 334682 700352
rect 397454 700340 397460 700352
rect 397512 700340 397518 700392
rect 480898 700340 480904 700392
rect 480956 700380 480962 700392
rect 494790 700380 494796 700392
rect 480956 700352 494796 700380
rect 480956 700340 480962 700352
rect 494790 700340 494796 700352
rect 494848 700340 494854 700392
rect 39850 700272 39856 700324
rect 39908 700312 39914 700324
rect 89162 700312 89168 700324
rect 39908 700284 89168 700312
rect 39908 700272 39914 700284
rect 89162 700272 89168 700284
rect 89220 700272 89226 700324
rect 137830 700272 137836 700324
rect 137888 700312 137894 700324
rect 176654 700312 176660 700324
rect 137888 700284 176660 700312
rect 137888 700272 137894 700284
rect 176654 700272 176660 700284
rect 176712 700272 176718 700324
rect 262858 700272 262864 700324
rect 262916 700312 262922 700324
rect 413646 700312 413652 700324
rect 262916 700284 413652 700312
rect 262916 700272 262922 700284
rect 413646 700272 413652 700284
rect 413704 700272 413710 700324
rect 479518 700272 479524 700324
rect 479576 700312 479582 700324
rect 559650 700312 559656 700324
rect 479576 700284 559656 700312
rect 479576 700272 479582 700284
rect 559650 700272 559656 700284
rect 559708 700272 559714 700324
rect 24302 699660 24308 699712
rect 24360 699700 24366 699712
rect 24762 699700 24768 699712
rect 24360 699672 24768 699700
rect 24360 699660 24366 699672
rect 24762 699660 24768 699672
rect 24820 699660 24826 699712
rect 39758 699660 39764 699712
rect 39816 699700 39822 699712
rect 40494 699700 40500 699712
rect 39816 699672 40500 699700
rect 39816 699660 39822 699672
rect 40494 699660 40500 699672
rect 40552 699660 40558 699712
rect 71774 699660 71780 699712
rect 71832 699700 71838 699712
rect 72970 699700 72976 699712
rect 71832 699672 72976 699700
rect 71832 699660 71838 699672
rect 72970 699660 72976 699672
rect 73028 699660 73034 699712
rect 266354 697552 266360 697604
rect 266412 697592 266418 697604
rect 267642 697592 267648 697604
rect 266412 697564 267648 697592
rect 266412 697552 266418 697564
rect 267642 697552 267648 697564
rect 267700 697552 267706 697604
rect 191098 696940 191104 696992
rect 191156 696980 191162 696992
rect 580166 696980 580172 696992
rect 191156 696952 580172 696980
rect 191156 696940 191162 696952
rect 580166 696940 580172 696952
rect 580224 696940 580230 696992
rect 2774 683612 2780 683664
rect 2832 683652 2838 683664
rect 6178 683652 6184 683664
rect 2832 683624 6184 683652
rect 2832 683612 2838 683624
rect 6178 683612 6184 683624
rect 6236 683612 6242 683664
rect 207658 683136 207664 683188
rect 207716 683176 207722 683188
rect 580166 683176 580172 683188
rect 207716 683148 580172 683176
rect 207716 683136 207722 683148
rect 580166 683136 580172 683148
rect 580224 683136 580230 683188
rect 182818 670692 182824 670744
rect 182876 670732 182882 670744
rect 580166 670732 580172 670744
rect 182876 670704 580172 670732
rect 182876 670692 182882 670704
rect 580166 670692 580172 670704
rect 580224 670692 580230 670744
rect 3510 656888 3516 656940
rect 3568 656928 3574 656940
rect 15838 656928 15844 656940
rect 3568 656900 15844 656928
rect 3568 656888 3574 656900
rect 15838 656888 15844 656900
rect 15896 656888 15902 656940
rect 189718 643084 189724 643136
rect 189776 643124 189782 643136
rect 580166 643124 580172 643136
rect 189776 643096 580172 643124
rect 189776 643084 189782 643096
rect 580166 643084 580172 643096
rect 580224 643084 580230 643136
rect 3510 632068 3516 632120
rect 3568 632108 3574 632120
rect 35158 632108 35164 632120
rect 3568 632080 35164 632108
rect 3568 632068 3574 632080
rect 35158 632068 35164 632080
rect 35216 632068 35222 632120
rect 180058 616836 180064 616888
rect 180116 616876 180122 616888
rect 580166 616876 580172 616888
rect 180116 616848 580172 616876
rect 180116 616836 180122 616848
rect 580166 616836 580172 616848
rect 580224 616836 580230 616888
rect 3326 605820 3332 605872
rect 3384 605860 3390 605872
rect 17218 605860 17224 605872
rect 3384 605832 17224 605860
rect 3384 605820 3390 605832
rect 17218 605820 17224 605832
rect 17276 605820 17282 605872
rect 258718 590656 258724 590708
rect 258776 590696 258782 590708
rect 580166 590696 580172 590708
rect 258776 590668 580172 590696
rect 258776 590656 258782 590668
rect 580166 590656 580172 590668
rect 580224 590656 580230 590708
rect 3326 579640 3332 579692
rect 3384 579680 3390 579692
rect 31018 579680 31024 579692
rect 3384 579652 31024 579680
rect 3384 579640 3390 579652
rect 31018 579640 31024 579652
rect 31076 579640 31082 579692
rect 204898 576852 204904 576904
rect 204956 576892 204962 576904
rect 580166 576892 580172 576904
rect 204956 576864 580172 576892
rect 204956 576852 204962 576864
rect 580166 576852 580172 576864
rect 580224 576852 580230 576904
rect 545758 563048 545764 563100
rect 545816 563088 545822 563100
rect 580166 563088 580172 563100
rect 545816 563060 580172 563088
rect 545816 563048 545822 563060
rect 580166 563048 580172 563060
rect 580224 563048 580230 563100
rect 3326 553392 3332 553444
rect 3384 553432 3390 553444
rect 28258 553432 28264 553444
rect 3384 553404 28264 553432
rect 3384 553392 3390 553404
rect 28258 553392 28264 553404
rect 28316 553392 28322 553444
rect 186958 536800 186964 536852
rect 187016 536840 187022 536852
rect 579890 536840 579896 536852
rect 187016 536812 579896 536840
rect 187016 536800 187022 536812
rect 579890 536800 579896 536812
rect 579948 536800 579954 536852
rect 3326 527144 3332 527196
rect 3384 527184 3390 527196
rect 10318 527184 10324 527196
rect 3384 527156 10324 527184
rect 3384 527144 3390 527156
rect 10318 527144 10324 527156
rect 10376 527144 10382 527196
rect 196618 524424 196624 524476
rect 196676 524464 196682 524476
rect 580166 524464 580172 524476
rect 196676 524436 580172 524464
rect 196676 524424 196682 524436
rect 580166 524424 580172 524436
rect 580224 524424 580230 524476
rect 3326 514768 3332 514820
rect 3384 514808 3390 514820
rect 32398 514808 32404 514820
rect 3384 514780 32404 514808
rect 3384 514768 3390 514780
rect 32398 514768 32404 514780
rect 32456 514768 32462 514820
rect 255958 510620 255964 510672
rect 256016 510660 256022 510672
rect 580166 510660 580172 510672
rect 256016 510632 580172 510660
rect 256016 510620 256022 510632
rect 580166 510620 580172 510632
rect 580224 510620 580230 510672
rect 2866 500964 2872 501016
rect 2924 501004 2930 501016
rect 33778 501004 33784 501016
rect 2924 500976 33784 501004
rect 2924 500964 2930 500976
rect 33778 500964 33784 500976
rect 33836 500964 33842 501016
rect 185578 484372 185584 484424
rect 185636 484412 185642 484424
rect 580166 484412 580172 484424
rect 185636 484384 580172 484412
rect 185636 484372 185642 484384
rect 580166 484372 580172 484384
rect 580224 484372 580230 484424
rect 3326 474716 3332 474768
rect 3384 474756 3390 474768
rect 13078 474756 13084 474768
rect 3384 474728 13084 474756
rect 3384 474716 3390 474728
rect 13078 474716 13084 474728
rect 13136 474716 13142 474768
rect 153194 473968 153200 474020
rect 153252 474008 153258 474020
rect 176746 474008 176752 474020
rect 153252 473980 176752 474008
rect 153252 473968 153258 473980
rect 176746 473968 176752 473980
rect 176804 473968 176810 474020
rect 3326 462340 3332 462392
rect 3384 462380 3390 462392
rect 21358 462380 21364 462392
rect 3384 462352 21364 462380
rect 3384 462340 3390 462352
rect 21358 462340 21364 462352
rect 21416 462340 21422 462392
rect 178678 456764 178684 456816
rect 178736 456804 178742 456816
rect 580166 456804 580172 456816
rect 178736 456776 580172 456804
rect 178736 456764 178742 456776
rect 580166 456764 580172 456776
rect 580224 456764 580230 456816
rect 3326 448536 3332 448588
rect 3384 448576 3390 448588
rect 19978 448576 19984 448588
rect 3384 448548 19984 448576
rect 3384 448536 3390 448548
rect 19978 448536 19984 448548
rect 20036 448536 20042 448588
rect 39666 425688 39672 425740
rect 39724 425728 39730 425740
rect 71774 425728 71780 425740
rect 39724 425700 71780 425728
rect 39724 425688 39730 425700
rect 71774 425688 71780 425700
rect 71832 425688 71838 425740
rect 106182 425688 106188 425740
rect 106240 425728 106246 425740
rect 176838 425728 176844 425740
rect 106240 425700 176844 425728
rect 106240 425688 106246 425700
rect 176838 425688 176844 425700
rect 176896 425688 176902 425740
rect 3142 422288 3148 422340
rect 3200 422328 3206 422340
rect 25498 422328 25504 422340
rect 3200 422300 25504 422328
rect 3200 422288 3206 422300
rect 25498 422288 25504 422300
rect 25556 422288 25562 422340
rect 486418 418140 486424 418192
rect 486476 418180 486482 418192
rect 580166 418180 580172 418192
rect 486476 418152 580172 418180
rect 486476 418140 486482 418152
rect 580166 418140 580172 418152
rect 580224 418140 580230 418192
rect 483658 404336 483664 404388
rect 483716 404376 483722 404388
rect 580166 404376 580172 404388
rect 483716 404348 580172 404376
rect 483716 404336 483722 404348
rect 580166 404336 580172 404348
rect 580224 404336 580230 404388
rect 3326 397468 3332 397520
rect 3384 397508 3390 397520
rect 21450 397508 21456 397520
rect 3384 397480 21456 397508
rect 3384 397468 3390 397480
rect 21450 397468 21456 397480
rect 21508 397468 21514 397520
rect 261478 376728 261484 376780
rect 261536 376768 261542 376780
rect 337654 376768 337660 376780
rect 261536 376740 337660 376768
rect 261536 376728 261542 376740
rect 337654 376728 337660 376740
rect 337712 376728 337718 376780
rect 254578 375368 254584 375420
rect 254636 375408 254642 375420
rect 337746 375408 337752 375420
rect 254636 375380 337752 375408
rect 254636 375368 254642 375380
rect 337746 375368 337752 375380
rect 337804 375368 337810 375420
rect 251818 372648 251824 372700
rect 251876 372688 251882 372700
rect 337470 372688 337476 372700
rect 251876 372660 337476 372688
rect 251876 372648 251882 372660
rect 337470 372648 337476 372660
rect 337528 372648 337534 372700
rect 198642 372580 198648 372632
rect 198700 372620 198706 372632
rect 337654 372620 337660 372632
rect 198700 372592 337660 372620
rect 198700 372580 198706 372592
rect 337654 372580 337660 372592
rect 337712 372580 337718 372632
rect 3326 371220 3332 371272
rect 3384 371260 3390 371272
rect 14458 371260 14464 371272
rect 3384 371232 14464 371260
rect 3384 371220 3390 371232
rect 14458 371220 14464 371232
rect 14516 371220 14522 371272
rect 250438 369928 250444 369980
rect 250496 369968 250502 369980
rect 337746 369968 337752 369980
rect 250496 369940 337752 369968
rect 250496 369928 250502 369940
rect 337746 369928 337752 369940
rect 337804 369928 337810 369980
rect 193122 369860 193128 369912
rect 193180 369900 193186 369912
rect 337470 369900 337476 369912
rect 193180 369872 337476 369900
rect 193180 369860 193186 369872
rect 337470 369860 337476 369872
rect 337528 369860 337534 369912
rect 249058 367072 249064 367124
rect 249116 367112 249122 367124
rect 337470 367112 337476 367124
rect 249116 367084 337476 367112
rect 249116 367072 249122 367084
rect 337470 367072 337476 367084
rect 337528 367072 337534 367124
rect 485038 364352 485044 364404
rect 485096 364392 485102 364404
rect 580166 364392 580172 364404
rect 485096 364364 580172 364392
rect 485096 364352 485102 364364
rect 580166 364352 580172 364364
rect 580224 364352 580230 364404
rect 482278 351908 482284 351960
rect 482336 351948 482342 351960
rect 580166 351948 580172 351960
rect 482336 351920 580172 351948
rect 482336 351908 482342 351920
rect 580166 351908 580172 351920
rect 580224 351908 580230 351960
rect 184842 349120 184848 349172
rect 184900 349160 184906 349172
rect 337286 349160 337292 349172
rect 184900 349132 337292 349160
rect 184900 349120 184906 349132
rect 337286 349120 337292 349132
rect 337344 349120 337350 349172
rect 33042 347828 33048 347880
rect 33100 347868 33106 347880
rect 37826 347868 37832 347880
rect 33100 347840 37832 347868
rect 33100 347828 33106 347840
rect 37826 347828 37832 347840
rect 37884 347828 37890 347880
rect 3050 345040 3056 345092
rect 3108 345080 3114 345092
rect 32490 345080 32496 345092
rect 3108 345052 32496 345080
rect 3108 345040 3114 345052
rect 32490 345040 32496 345052
rect 32548 345040 32554 345092
rect 38102 339396 38108 339448
rect 38160 339436 38166 339448
rect 131758 339436 131764 339448
rect 38160 339408 131764 339436
rect 38160 339396 38166 339408
rect 131758 339396 131764 339408
rect 131816 339396 131822 339448
rect 38286 339328 38292 339380
rect 38344 339368 38350 339380
rect 153838 339368 153844 339380
rect 38344 339340 153844 339368
rect 38344 339328 38350 339340
rect 153838 339328 153844 339340
rect 153896 339328 153902 339380
rect 3418 339260 3424 339312
rect 3476 339300 3482 339312
rect 132494 339300 132500 339312
rect 3476 339272 132500 339300
rect 3476 339260 3482 339272
rect 132494 339260 132500 339272
rect 132552 339260 132558 339312
rect 3510 339192 3516 339244
rect 3568 339232 3574 339244
rect 136634 339232 136640 339244
rect 3568 339204 136640 339232
rect 3568 339192 3574 339204
rect 136634 339192 136640 339204
rect 136692 339192 136698 339244
rect 3602 339124 3608 339176
rect 3660 339164 3666 339176
rect 140774 339164 140780 339176
rect 3660 339136 140780 339164
rect 3660 339124 3666 339136
rect 140774 339124 140780 339136
rect 140832 339124 140838 339176
rect 3786 339056 3792 339108
rect 3844 339096 3850 339108
rect 155954 339096 155960 339108
rect 3844 339068 155960 339096
rect 3844 339056 3850 339068
rect 155954 339056 155960 339068
rect 156012 339056 156018 339108
rect 38838 338988 38844 339040
rect 38896 339028 38902 339040
rect 193214 339028 193220 339040
rect 38896 339000 193220 339028
rect 38896 338988 38902 339000
rect 193214 338988 193220 339000
rect 193272 338988 193278 339040
rect 92290 338920 92296 338972
rect 92348 338960 92354 338972
rect 580258 338960 580264 338972
rect 92348 338932 580264 338960
rect 92348 338920 92354 338932
rect 580258 338920 580264 338932
rect 580316 338920 580322 338972
rect 81342 338852 81348 338904
rect 81400 338892 81406 338904
rect 580350 338892 580356 338904
rect 81400 338864 580356 338892
rect 81400 338852 81406 338864
rect 580350 338852 580356 338864
rect 580408 338852 580414 338904
rect 75822 338784 75828 338836
rect 75880 338824 75886 338836
rect 580442 338824 580448 338836
rect 75880 338796 580448 338824
rect 75880 338784 75886 338796
rect 580442 338784 580448 338796
rect 580500 338784 580506 338836
rect 73062 338716 73068 338768
rect 73120 338756 73126 338768
rect 580534 338756 580540 338768
rect 73120 338728 580540 338756
rect 73120 338716 73126 338728
rect 580534 338716 580540 338728
rect 580592 338716 580598 338768
rect 39758 338648 39764 338700
rect 39816 338688 39822 338700
rect 126974 338688 126980 338700
rect 39816 338660 126980 338688
rect 39816 338648 39822 338660
rect 126974 338648 126980 338660
rect 127032 338648 127038 338700
rect 38562 338036 38568 338088
rect 38620 338076 38626 338088
rect 337378 338076 337384 338088
rect 38620 338048 337384 338076
rect 38620 338036 38626 338048
rect 337378 338036 337384 338048
rect 337436 338036 337442 338088
rect 48958 337968 48964 338020
rect 49016 338008 49022 338020
rect 368474 338008 368480 338020
rect 49016 337980 368480 338008
rect 49016 337968 49022 337980
rect 368474 337968 368480 337980
rect 368532 337968 368538 338020
rect 40494 337900 40500 337952
rect 40552 337940 40558 337952
rect 356054 337940 356060 337952
rect 40552 337912 356060 337940
rect 40552 337900 40558 337912
rect 356054 337900 356060 337912
rect 356112 337900 356118 337952
rect 56502 337832 56508 337884
rect 56560 337872 56566 337884
rect 236638 337872 236644 337884
rect 56560 337844 236644 337872
rect 56560 337832 56566 337844
rect 236638 337832 236644 337844
rect 236696 337832 236702 337884
rect 43438 337764 43444 337816
rect 43496 337804 43502 337816
rect 394694 337804 394700 337816
rect 43496 337776 394700 337804
rect 43496 337764 43502 337776
rect 394694 337764 394700 337776
rect 394752 337764 394758 337816
rect 99282 337696 99288 337748
rect 99340 337736 99346 337748
rect 226978 337736 226984 337748
rect 99340 337708 226984 337736
rect 99340 337696 99346 337708
rect 226978 337696 226984 337708
rect 227036 337696 227042 337748
rect 95142 337628 95148 337680
rect 95200 337668 95206 337680
rect 225598 337668 225604 337680
rect 95200 337640 225604 337668
rect 95200 337628 95206 337640
rect 225598 337628 225604 337640
rect 225656 337628 225662 337680
rect 385678 337628 385684 337680
rect 385736 337668 385742 337680
rect 387794 337668 387800 337680
rect 385736 337640 387800 337668
rect 385736 337628 385742 337640
rect 387794 337628 387800 337640
rect 387852 337628 387858 337680
rect 388438 337628 388444 337680
rect 388496 337668 388502 337680
rect 390554 337668 390560 337680
rect 388496 337640 390560 337668
rect 388496 337628 388502 337640
rect 390554 337628 390560 337640
rect 390612 337628 390618 337680
rect 91002 337560 91008 337612
rect 91060 337600 91066 337612
rect 239398 337600 239404 337612
rect 91060 337572 239404 337600
rect 91060 337560 91066 337572
rect 239398 337560 239404 337572
rect 239456 337560 239462 337612
rect 387058 337560 387064 337612
rect 387116 337600 387122 337612
rect 389174 337600 389180 337612
rect 387116 337572 389180 337600
rect 387116 337560 387122 337572
rect 389174 337560 389180 337572
rect 389232 337560 389238 337612
rect 78582 337492 78588 337544
rect 78640 337532 78646 337544
rect 239582 337532 239588 337544
rect 78640 337504 239588 337532
rect 78640 337492 78646 337504
rect 239582 337492 239588 337504
rect 239640 337492 239646 337544
rect 77202 337424 77208 337476
rect 77260 337464 77266 337476
rect 239490 337464 239496 337476
rect 77260 337436 239496 337464
rect 77260 337424 77266 337436
rect 239490 337424 239496 337436
rect 239548 337424 239554 337476
rect 57882 337356 57888 337408
rect 57940 337396 57946 337408
rect 221458 337396 221464 337408
rect 57940 337368 221464 337396
rect 57940 337356 57946 337368
rect 221458 337356 221464 337368
rect 221516 337356 221522 337408
rect 359458 337356 359464 337408
rect 359516 337396 359522 337408
rect 378134 337396 378140 337408
rect 359516 337368 378140 337396
rect 359516 337356 359522 337368
rect 378134 337356 378140 337368
rect 378192 337356 378198 337408
rect 216582 337288 216588 337340
rect 216640 337328 216646 337340
rect 382274 337328 382280 337340
rect 216640 337300 382280 337328
rect 216640 337288 216646 337300
rect 382274 337288 382280 337300
rect 382332 337288 382338 337340
rect 382918 337288 382924 337340
rect 382976 337328 382982 337340
rect 390554 337328 390560 337340
rect 382976 337300 390560 337328
rect 382976 337288 382982 337300
rect 390554 337288 390560 337300
rect 390612 337288 390618 337340
rect 391290 337288 391296 337340
rect 391348 337328 391354 337340
rect 397454 337328 397460 337340
rect 391348 337300 397460 337328
rect 391348 337288 391354 337300
rect 397454 337288 397460 337300
rect 397512 337288 397518 337340
rect 40402 337220 40408 337272
rect 40460 337260 40466 337272
rect 59446 337260 59452 337272
rect 40460 337232 59452 337260
rect 40460 337220 40466 337232
rect 59446 337220 59452 337232
rect 59504 337220 59510 337272
rect 72970 337220 72976 337272
rect 73028 337260 73034 337272
rect 239674 337260 239680 337272
rect 73028 337232 239680 337260
rect 73028 337220 73034 337232
rect 239674 337220 239680 337232
rect 239732 337220 239738 337272
rect 240042 337220 240048 337272
rect 240100 337260 240106 337272
rect 398834 337260 398840 337272
rect 240100 337232 398840 337260
rect 240100 337220 240106 337232
rect 398834 337220 398840 337232
rect 398892 337220 398898 337272
rect 39390 337152 39396 337204
rect 39448 337192 39454 337204
rect 59354 337192 59360 337204
rect 39448 337164 59360 337192
rect 39448 337152 39454 337164
rect 59354 337152 59360 337164
rect 59412 337152 59418 337204
rect 203518 337152 203524 337204
rect 203576 337192 203582 337204
rect 371234 337192 371240 337204
rect 203576 337164 371240 337192
rect 203576 337152 203582 337164
rect 371234 337152 371240 337164
rect 371292 337152 371298 337204
rect 373258 337152 373264 337204
rect 373316 337192 373322 337204
rect 445754 337192 445760 337204
rect 373316 337164 445760 337192
rect 373316 337152 373322 337164
rect 445754 337152 445760 337164
rect 445812 337152 445818 337204
rect 234522 337084 234528 337136
rect 234580 337124 234586 337136
rect 396074 337124 396080 337136
rect 234580 337096 396080 337124
rect 234580 337084 234586 337096
rect 396074 337084 396080 337096
rect 396132 337084 396138 337136
rect 355318 337016 355324 337068
rect 355376 337056 355382 337068
rect 375374 337056 375380 337068
rect 355376 337028 375380 337056
rect 355376 337016 355382 337028
rect 375374 337016 375380 337028
rect 375432 337016 375438 337068
rect 377398 337016 377404 337068
rect 377456 337056 377462 337068
rect 391934 337056 391940 337068
rect 377456 337028 391940 337056
rect 377456 337016 377462 337028
rect 391934 337016 391940 337028
rect 391992 337016 391998 337068
rect 42058 336948 42064 337000
rect 42116 336988 42122 337000
rect 361574 336988 361580 337000
rect 42116 336960 361580 336988
rect 42116 336948 42122 336960
rect 361574 336948 361580 336960
rect 361632 336948 361638 337000
rect 370498 336948 370504 337000
rect 370556 336988 370562 337000
rect 437474 336988 437480 337000
rect 370556 336960 437480 336988
rect 370556 336948 370562 336960
rect 437474 336948 437480 336960
rect 437532 336948 437538 337000
rect 367738 336880 367744 336932
rect 367796 336920 367802 336932
rect 434714 336920 434720 336932
rect 367796 336892 434720 336920
rect 367796 336880 367802 336892
rect 434714 336880 434720 336892
rect 434772 336880 434778 336932
rect 50338 336812 50344 336864
rect 50396 336852 50402 336864
rect 369854 336852 369860 336864
rect 50396 336824 369860 336852
rect 50396 336812 50402 336824
rect 369854 336812 369860 336824
rect 369912 336812 369918 336864
rect 93578 336744 93584 336796
rect 93636 336784 93642 336796
rect 100018 336784 100024 336796
rect 93636 336756 100024 336784
rect 93636 336744 93642 336756
rect 100018 336744 100024 336756
rect 100076 336744 100082 336796
rect 391198 336744 391204 336796
rect 391256 336784 391262 336796
rect 393866 336784 393872 336796
rect 391256 336756 393872 336784
rect 391256 336744 391262 336756
rect 393866 336744 393872 336756
rect 393924 336744 393930 336796
rect 420178 336744 420184 336796
rect 420236 336784 420242 336796
rect 422662 336784 422668 336796
rect 420236 336756 422668 336784
rect 420236 336744 420242 336756
rect 422662 336744 422668 336756
rect 422720 336744 422726 336796
rect 119982 336540 119988 336592
rect 120040 336580 120046 336592
rect 178034 336580 178040 336592
rect 120040 336552 178040 336580
rect 120040 336540 120046 336552
rect 178034 336540 178040 336552
rect 178092 336540 178098 336592
rect 99282 336472 99288 336524
rect 99340 336512 99346 336524
rect 171778 336512 171784 336524
rect 99340 336484 171784 336512
rect 99340 336472 99346 336484
rect 171778 336472 171784 336484
rect 171836 336472 171842 336524
rect 96522 336404 96528 336456
rect 96580 336444 96586 336456
rect 173158 336444 173164 336456
rect 96580 336416 173164 336444
rect 96580 336404 96586 336416
rect 173158 336404 173164 336416
rect 173216 336404 173222 336456
rect 131022 336336 131028 336388
rect 131080 336376 131086 336388
rect 213178 336376 213184 336388
rect 131080 336348 213184 336376
rect 131080 336336 131086 336348
rect 213178 336336 213184 336348
rect 213236 336336 213242 336388
rect 81250 336268 81256 336320
rect 81308 336308 81314 336320
rect 177298 336308 177304 336320
rect 81308 336280 177304 336308
rect 81308 336268 81314 336280
rect 177298 336268 177304 336280
rect 177356 336268 177362 336320
rect 117222 336200 117228 336252
rect 117280 336240 117286 336252
rect 214558 336240 214564 336252
rect 117280 336212 214564 336240
rect 117280 336200 117286 336212
rect 214558 336200 214564 336212
rect 214616 336200 214622 336252
rect 229738 336200 229744 336252
rect 229796 336240 229802 336252
rect 385126 336240 385132 336252
rect 229796 336212 385132 336240
rect 229796 336200 229802 336212
rect 385126 336200 385132 336212
rect 385184 336200 385190 336252
rect 77202 336132 77208 336184
rect 77260 336172 77266 336184
rect 242894 336172 242900 336184
rect 77260 336144 242900 336172
rect 77260 336132 77266 336144
rect 242894 336132 242900 336144
rect 242952 336132 242958 336184
rect 247678 336132 247684 336184
rect 247736 336172 247742 336184
rect 369946 336172 369952 336184
rect 247736 336144 369952 336172
rect 247736 336132 247742 336144
rect 369946 336132 369952 336144
rect 370004 336132 370010 336184
rect 32398 336064 32404 336116
rect 32456 336104 32462 336116
rect 143534 336104 143540 336116
rect 32456 336076 143540 336104
rect 32456 336064 32462 336076
rect 143534 336064 143540 336076
rect 143592 336064 143598 336116
rect 209682 336064 209688 336116
rect 209740 336104 209746 336116
rect 400214 336104 400220 336116
rect 209740 336076 400220 336104
rect 209740 336064 209746 336076
rect 400214 336064 400220 336076
rect 400272 336064 400278 336116
rect 34422 335996 34428 336048
rect 34480 336036 34486 336048
rect 382274 336036 382280 336048
rect 34480 336008 382280 336036
rect 34480 335996 34486 336008
rect 382274 335996 382280 336008
rect 382332 335996 382338 336048
rect 81066 334908 81072 334960
rect 81124 334948 81130 334960
rect 200758 334948 200764 334960
rect 81124 334920 200764 334948
rect 81124 334908 81130 334920
rect 200758 334908 200764 334920
rect 200816 334908 200822 334960
rect 74902 334840 74908 334892
rect 74960 334880 74966 334892
rect 195238 334880 195244 334892
rect 74960 334852 195244 334880
rect 74960 334840 74966 334852
rect 195238 334840 195244 334852
rect 195296 334840 195302 334892
rect 76282 334772 76288 334824
rect 76340 334812 76346 334824
rect 243078 334812 243084 334824
rect 76340 334784 243084 334812
rect 76340 334772 76346 334784
rect 243078 334772 243084 334784
rect 243136 334772 243142 334824
rect 31386 334704 31392 334756
rect 31444 334744 31450 334756
rect 386598 334744 386604 334756
rect 31444 334716 386604 334744
rect 31444 334704 31450 334716
rect 386598 334704 386604 334716
rect 386656 334704 386662 334756
rect 35710 334636 35716 334688
rect 35768 334676 35774 334688
rect 396166 334676 396172 334688
rect 35768 334648 396172 334676
rect 35768 334636 35774 334648
rect 396166 334636 396172 334648
rect 396224 334636 396230 334688
rect 34330 334568 34336 334620
rect 34388 334608 34394 334620
rect 407114 334608 407120 334620
rect 34388 334580 407120 334608
rect 34388 334568 34394 334580
rect 407114 334568 407120 334580
rect 407172 334568 407178 334620
rect 85298 333548 85304 333600
rect 85356 333588 85362 333600
rect 162118 333588 162124 333600
rect 85356 333560 162124 333588
rect 85356 333548 85362 333560
rect 162118 333548 162124 333560
rect 162176 333548 162182 333600
rect 86402 333480 86408 333532
rect 86460 333520 86466 333532
rect 169018 333520 169024 333532
rect 86460 333492 169024 333520
rect 86460 333480 86466 333492
rect 169018 333480 169024 333492
rect 169076 333480 169082 333532
rect 90634 333412 90640 333464
rect 90692 333452 90698 333464
rect 220078 333452 220084 333464
rect 90692 333424 220084 333452
rect 90692 333412 90698 333424
rect 220078 333412 220084 333424
rect 220136 333412 220142 333464
rect 38654 333344 38660 333396
rect 38712 333384 38718 333396
rect 189074 333384 189080 333396
rect 38712 333356 189080 333384
rect 38712 333344 38718 333356
rect 189074 333344 189080 333356
rect 189132 333344 189138 333396
rect 83550 333276 83556 333328
rect 83608 333316 83614 333328
rect 244458 333316 244464 333328
rect 83608 333288 244464 333316
rect 83608 333276 83614 333288
rect 244458 333276 244464 333288
rect 244516 333276 244522 333328
rect 30282 333208 30288 333260
rect 30340 333248 30346 333260
rect 360194 333248 360200 333260
rect 30340 333220 360200 333248
rect 30340 333208 30346 333220
rect 360194 333208 360200 333220
rect 360252 333208 360258 333260
rect 38654 324912 38660 324964
rect 38712 324952 38718 324964
rect 67634 324952 67640 324964
rect 38712 324924 67640 324952
rect 38712 324912 38718 324924
rect 67634 324912 67640 324924
rect 67692 324912 67698 324964
rect 68830 324300 68836 324352
rect 68888 324340 68894 324352
rect 580166 324340 580172 324352
rect 68888 324312 580172 324340
rect 68888 324300 68894 324312
rect 580166 324300 580172 324312
rect 580224 324300 580230 324352
rect 3418 318792 3424 318844
rect 3476 318832 3482 318844
rect 156046 318832 156052 318844
rect 3476 318804 156052 318832
rect 3476 318792 3482 318804
rect 156046 318792 156052 318804
rect 156104 318792 156110 318844
rect 70302 311856 70308 311908
rect 70360 311896 70366 311908
rect 580166 311896 580172 311908
rect 70360 311868 580172 311896
rect 70360 311856 70366 311868
rect 580166 311856 580172 311868
rect 580224 311856 580230 311908
rect 21450 311108 21456 311160
rect 21508 311148 21514 311160
rect 150434 311148 150440 311160
rect 21508 311120 150440 311148
rect 21508 311108 21514 311120
rect 150434 311108 150440 311120
rect 150492 311108 150498 311160
rect 3418 304988 3424 305040
rect 3476 305028 3482 305040
rect 158714 305028 158720 305040
rect 3476 305000 158720 305028
rect 3476 304988 3482 305000
rect 158714 304988 158720 305000
rect 158772 304988 158778 305040
rect 67542 298120 67548 298172
rect 67600 298160 67606 298172
rect 580166 298160 580172 298172
rect 67600 298132 580172 298160
rect 67600 298120 67606 298132
rect 580166 298120 580172 298132
rect 580224 298120 580230 298172
rect 32858 297372 32864 297424
rect 32916 297412 32922 297424
rect 387886 297412 387892 297424
rect 32916 297384 387892 297412
rect 32916 297372 32922 297384
rect 387886 297372 387892 297384
rect 387944 297372 387950 297424
rect 3418 292544 3424 292596
rect 3476 292584 3482 292596
rect 157334 292584 157340 292596
rect 3476 292556 157340 292584
rect 3476 292544 3482 292556
rect 157334 292544 157340 292556
rect 157392 292544 157398 292596
rect 19978 290436 19984 290488
rect 20036 290476 20042 290488
rect 146294 290476 146300 290488
rect 20036 290448 146300 290476
rect 20036 290436 20042 290448
rect 146294 290436 146300 290448
rect 146352 290436 146358 290488
rect 28258 282140 28264 282192
rect 28316 282180 28322 282192
rect 139394 282180 139400 282192
rect 28316 282152 139400 282180
rect 28316 282140 28322 282152
rect 139394 282140 139400 282152
rect 139452 282140 139458 282192
rect 25498 280780 25504 280832
rect 25556 280820 25562 280832
rect 149054 280820 149060 280832
rect 25556 280792 149060 280820
rect 25556 280780 25562 280792
rect 149054 280780 149060 280792
rect 149112 280780 149118 280832
rect 38746 277992 38752 278044
rect 38804 278032 38810 278044
rect 241514 278032 241520 278044
rect 38804 278004 241520 278032
rect 38804 277992 38810 278004
rect 241514 277992 241520 278004
rect 241572 277992 241578 278044
rect 31662 275272 31668 275324
rect 31720 275312 31726 275324
rect 364334 275312 364340 275324
rect 31720 275284 364340 275312
rect 31720 275272 31726 275284
rect 364334 275272 364340 275284
rect 364392 275272 364398 275324
rect 97902 273912 97908 273964
rect 97960 273952 97966 273964
rect 232498 273952 232504 273964
rect 97960 273924 232504 273952
rect 97960 273912 97966 273924
rect 232498 273912 232504 273924
rect 232556 273912 232562 273964
rect 64690 271872 64696 271924
rect 64748 271912 64754 271924
rect 579798 271912 579804 271924
rect 64748 271884 579804 271912
rect 64748 271872 64754 271884
rect 579798 271872 579804 271884
rect 579856 271872 579862 271924
rect 100018 271124 100024 271176
rect 100076 271164 100082 271176
rect 230474 271164 230480 271176
rect 100076 271136 230480 271164
rect 100076 271124 100082 271136
rect 230474 271124 230480 271136
rect 230532 271124 230538 271176
rect 79962 269764 79968 269816
rect 80020 269804 80026 269816
rect 244642 269804 244648 269816
rect 80020 269776 244648 269804
rect 80020 269764 80026 269776
rect 244642 269764 244648 269776
rect 244700 269764 244706 269816
rect 88150 268336 88156 268388
rect 88208 268376 88214 268388
rect 167638 268376 167644 268388
rect 88208 268348 167644 268376
rect 88208 268336 88214 268348
rect 167638 268336 167644 268348
rect 167696 268336 167702 268388
rect 3050 266364 3056 266416
rect 3108 266404 3114 266416
rect 160554 266404 160560 266416
rect 3108 266376 160560 266404
rect 3108 266364 3114 266376
rect 160554 266364 160560 266376
rect 160612 266364 160618 266416
rect 126882 265616 126888 265668
rect 126940 265656 126946 265668
rect 222838 265656 222844 265668
rect 126940 265628 222844 265656
rect 126940 265616 126946 265628
rect 222838 265616 222844 265628
rect 222896 265616 222902 265668
rect 107562 264256 107568 264308
rect 107620 264296 107626 264308
rect 262858 264296 262864 264308
rect 107620 264268 262864 264296
rect 107620 264256 107626 264268
rect 262858 264256 262864 264268
rect 262916 264256 262922 264308
rect 34238 264188 34244 264240
rect 34296 264228 34302 264240
rect 380986 264228 380992 264240
rect 34296 264200 380992 264228
rect 34296 264188 34302 264200
rect 380986 264188 380992 264200
rect 381044 264188 381050 264240
rect 85482 262828 85488 262880
rect 85540 262868 85546 262880
rect 196618 262868 196624 262880
rect 85540 262840 196624 262868
rect 85540 262828 85546 262840
rect 196618 262828 196624 262840
rect 196676 262828 196682 262880
rect 100018 261468 100024 261520
rect 100076 261508 100082 261520
rect 527174 261508 527180 261520
rect 100076 261480 527180 261508
rect 100076 261468 100082 261480
rect 527174 261468 527180 261480
rect 527232 261468 527238 261520
rect 32490 260176 32496 260228
rect 32548 260216 32554 260228
rect 154574 260216 154580 260228
rect 32548 260188 154580 260216
rect 32548 260176 32554 260188
rect 154574 260176 154580 260188
rect 154632 260176 154638 260228
rect 88150 260108 88156 260160
rect 88208 260148 88214 260160
rect 258718 260148 258724 260160
rect 88208 260120 258724 260148
rect 88208 260108 88214 260120
rect 258718 260108 258724 260120
rect 258776 260108 258782 260160
rect 66162 258068 66168 258120
rect 66220 258108 66226 258120
rect 580166 258108 580172 258120
rect 66220 258080 580172 258108
rect 66220 258068 66226 258080
rect 580166 258068 580172 258080
rect 580224 258068 580230 258120
rect 71682 257320 71688 257372
rect 71740 257360 71746 257372
rect 482278 257360 482284 257372
rect 71740 257332 482284 257360
rect 71740 257320 71746 257332
rect 482278 257320 482284 257332
rect 482336 257320 482342 257372
rect 36998 255960 37004 256012
rect 37056 256000 37062 256012
rect 92474 256000 92480 256012
rect 37056 255972 92480 256000
rect 37056 255960 37062 255972
rect 92474 255960 92480 255972
rect 92532 255960 92538 256012
rect 108758 255960 108764 256012
rect 108816 256000 108822 256012
rect 333238 256000 333244 256012
rect 108816 255972 333244 256000
rect 108816 255960 108822 255972
rect 333238 255960 333244 255972
rect 333296 255960 333302 256012
rect 78490 254600 78496 254652
rect 78548 254640 78554 254652
rect 244550 254640 244556 254652
rect 78548 254612 244556 254640
rect 78548 254600 78554 254612
rect 244550 254600 244556 254612
rect 244608 254600 244614 254652
rect 74350 254532 74356 254584
rect 74408 254572 74414 254584
rect 245654 254572 245660 254584
rect 74408 254544 245660 254572
rect 74408 254532 74414 254544
rect 245654 254532 245660 254544
rect 245712 254532 245718 254584
rect 3418 253920 3424 253972
rect 3476 253960 3482 253972
rect 163130 253960 163136 253972
rect 3476 253932 163136 253960
rect 3476 253920 3482 253932
rect 163130 253920 163136 253932
rect 163188 253920 163194 253972
rect 35802 253580 35808 253632
rect 35860 253620 35866 253632
rect 135254 253620 135260 253632
rect 35860 253592 135260 253620
rect 35860 253580 35866 253592
rect 135254 253580 135260 253592
rect 135312 253580 135318 253632
rect 118602 253512 118608 253564
rect 118660 253552 118666 253564
rect 220814 253552 220820 253564
rect 118660 253524 220820 253552
rect 118660 253512 118666 253524
rect 220814 253512 220820 253524
rect 220872 253512 220878 253564
rect 129642 253444 129648 253496
rect 129700 253484 129706 253496
rect 243446 253484 243452 253496
rect 129700 253456 243452 253484
rect 129700 253444 129706 253456
rect 243446 253444 243452 253456
rect 243504 253444 243510 253496
rect 21358 253376 21364 253428
rect 21416 253416 21422 253428
rect 148042 253416 148048 253428
rect 21416 253388 148048 253416
rect 21416 253376 21422 253388
rect 148042 253376 148048 253388
rect 148100 253376 148106 253428
rect 104710 253308 104716 253360
rect 104768 253348 104774 253360
rect 327718 253348 327724 253360
rect 104768 253320 327724 253348
rect 104768 253308 104774 253320
rect 327718 253308 327724 253320
rect 327776 253308 327782 253360
rect 31478 253240 31484 253292
rect 31536 253280 31542 253292
rect 367186 253280 367192 253292
rect 31536 253252 367192 253280
rect 31536 253240 31542 253252
rect 367186 253240 367192 253252
rect 367244 253240 367250 253292
rect 33962 253172 33968 253224
rect 34020 253212 34026 253224
rect 409874 253212 409880 253224
rect 34020 253184 409880 253212
rect 34020 253172 34026 253184
rect 409874 253172 409880 253184
rect 409932 253172 409938 253224
rect 117958 252356 117964 252408
rect 118016 252396 118022 252408
rect 201494 252396 201500 252408
rect 118016 252368 201500 252396
rect 118016 252356 118022 252368
rect 201494 252356 201500 252368
rect 201552 252356 201558 252408
rect 111610 252288 111616 252340
rect 111668 252328 111674 252340
rect 211798 252328 211804 252340
rect 111668 252300 211804 252328
rect 111668 252288 111674 252300
rect 211798 252288 211804 252300
rect 211856 252288 211862 252340
rect 17218 252220 17224 252272
rect 17276 252260 17282 252272
rect 135530 252260 135536 252272
rect 17276 252232 135536 252260
rect 17276 252220 17282 252232
rect 135530 252220 135536 252232
rect 135588 252220 135594 252272
rect 14458 252152 14464 252204
rect 14516 252192 14522 252204
rect 153194 252192 153200 252204
rect 14516 252164 153200 252192
rect 14516 252152 14522 252164
rect 153194 252152 153200 252164
rect 153252 252152 153258 252204
rect 35434 252084 35440 252136
rect 35492 252124 35498 252136
rect 113174 252124 113180 252136
rect 35492 252096 113180 252124
rect 35492 252084 35498 252096
rect 113174 252084 113180 252096
rect 113232 252084 113238 252136
rect 114462 252084 114468 252136
rect 114520 252124 114526 252136
rect 266354 252124 266360 252136
rect 114520 252096 266360 252124
rect 114520 252084 114526 252096
rect 266354 252084 266360 252096
rect 266412 252084 266418 252136
rect 74442 252016 74448 252068
rect 74500 252056 74506 252068
rect 243170 252056 243176 252068
rect 74500 252028 243176 252056
rect 74500 252016 74506 252028
rect 243170 252016 243176 252028
rect 243228 252016 243234 252068
rect 106090 251948 106096 252000
rect 106148 251988 106154 252000
rect 334618 251988 334624 252000
rect 106148 251960 334624 251988
rect 106148 251948 106154 251960
rect 334618 251948 334624 251960
rect 334676 251948 334682 252000
rect 32674 251880 32680 251932
rect 32732 251920 32738 251932
rect 383654 251920 383660 251932
rect 32732 251892 383660 251920
rect 32732 251880 32738 251892
rect 383654 251880 383660 251892
rect 383712 251880 383718 251932
rect 102042 251812 102048 251864
rect 102100 251852 102106 251864
rect 480898 251852 480904 251864
rect 102100 251824 480904 251852
rect 102100 251812 102106 251824
rect 480898 251812 480904 251824
rect 480956 251812 480962 251864
rect 109494 251064 109500 251116
rect 109552 251104 109558 251116
rect 193858 251104 193864 251116
rect 109552 251076 193864 251104
rect 109552 251064 109558 251076
rect 193858 251064 193864 251076
rect 193916 251064 193922 251116
rect 90726 250996 90732 251048
rect 90784 251036 90790 251048
rect 189718 251036 189724 251048
rect 90784 251008 189724 251036
rect 90784 250996 90790 251008
rect 189718 250996 189724 251008
rect 189776 250996 189782 251048
rect 37090 250928 37096 250980
rect 37148 250968 37154 250980
rect 142154 250968 142160 250980
rect 37148 250940 142160 250968
rect 37148 250928 37154 250940
rect 142154 250928 142160 250940
rect 142212 250928 142218 250980
rect 79410 250860 79416 250912
rect 79468 250900 79474 250912
rect 185578 250900 185584 250912
rect 79468 250872 185584 250900
rect 79468 250860 79474 250872
rect 185578 250860 185584 250872
rect 185636 250860 185642 250912
rect 15838 250792 15844 250844
rect 15896 250832 15902 250844
rect 132126 250832 132132 250844
rect 15896 250804 132132 250832
rect 15896 250792 15902 250804
rect 132126 250792 132132 250804
rect 132184 250792 132190 250844
rect 142062 250792 142068 250844
rect 142120 250832 142126 250844
rect 242986 250832 242992 250844
rect 142120 250804 242992 250832
rect 142120 250792 142126 250804
rect 242986 250792 242992 250804
rect 243044 250792 243050 250844
rect 10318 250724 10324 250776
rect 10376 250764 10382 250776
rect 142154 250764 142160 250776
rect 10376 250736 142160 250764
rect 10376 250724 10382 250736
rect 142154 250724 142160 250736
rect 142212 250724 142218 250776
rect 106182 250656 106188 250708
rect 106240 250696 106246 250708
rect 240502 250696 240508 250708
rect 106240 250668 240508 250696
rect 106240 250656 106246 250668
rect 240502 250656 240508 250668
rect 240560 250656 240566 250708
rect 81894 250588 81900 250640
rect 81952 250628 81958 250640
rect 255958 250628 255964 250640
rect 81952 250600 255964 250628
rect 81952 250588 81958 250600
rect 255958 250588 255964 250600
rect 256016 250588 256022 250640
rect 36906 250520 36912 250572
rect 36964 250560 36970 250572
rect 100754 250560 100760 250572
rect 36964 250532 100760 250560
rect 36964 250520 36970 250532
rect 100754 250520 100760 250532
rect 100812 250520 100818 250572
rect 101950 250520 101956 250572
rect 102008 250560 102014 250572
rect 330478 250560 330484 250572
rect 102008 250532 330484 250560
rect 102008 250520 102014 250532
rect 330478 250520 330484 250532
rect 330536 250520 330542 250572
rect 74442 250452 74448 250504
rect 74500 250492 74506 250504
rect 483658 250492 483664 250504
rect 74500 250464 483664 250492
rect 74500 250452 74506 250464
rect 483658 250452 483664 250464
rect 483716 250452 483722 250504
rect 93210 249704 93216 249756
rect 93268 249744 93274 249756
rect 182818 249744 182824 249756
rect 93268 249716 182824 249744
rect 93268 249704 93274 249716
rect 182818 249704 182824 249716
rect 182876 249704 182882 249756
rect 89438 249636 89444 249688
rect 89496 249676 89502 249688
rect 180058 249676 180064 249688
rect 89496 249648 180064 249676
rect 89496 249636 89502 249648
rect 180058 249636 180064 249648
rect 180116 249636 180122 249688
rect 36722 249568 36728 249620
rect 36780 249608 36786 249620
rect 122834 249608 122840 249620
rect 36780 249580 122840 249608
rect 36780 249568 36786 249580
rect 122834 249568 122840 249580
rect 122892 249568 122898 249620
rect 146202 249568 146208 249620
rect 146260 249608 146266 249620
rect 239766 249608 239772 249620
rect 146260 249580 239772 249608
rect 146260 249568 146266 249580
rect 239766 249568 239772 249580
rect 239824 249568 239830 249620
rect 94498 249500 94504 249552
rect 94556 249540 94562 249552
rect 191098 249540 191104 249552
rect 94556 249512 191104 249540
rect 94556 249500 94562 249512
rect 191098 249500 191104 249512
rect 191156 249500 191162 249552
rect 78214 249432 78220 249484
rect 78272 249472 78278 249484
rect 178678 249472 178684 249484
rect 78272 249444 178684 249472
rect 78272 249432 78278 249444
rect 178678 249432 178684 249444
rect 178736 249432 178742 249484
rect 83182 249364 83188 249416
rect 83240 249404 83246 249416
rect 186958 249404 186964 249416
rect 83240 249376 186964 249404
rect 83240 249364 83246 249376
rect 186958 249364 186964 249376
rect 187016 249364 187022 249416
rect 121362 249296 121368 249348
rect 121420 249336 121426 249348
rect 240134 249336 240140 249348
rect 121420 249308 240140 249336
rect 121420 249296 121426 249308
rect 240134 249296 240140 249308
rect 240192 249296 240198 249348
rect 104802 249228 104808 249280
rect 104860 249268 104866 249280
rect 240410 249268 240416 249280
rect 104860 249240 240416 249268
rect 104860 249228 104866 249240
rect 240410 249228 240416 249240
rect 240468 249228 240474 249280
rect 6178 249160 6184 249212
rect 6236 249200 6242 249212
rect 130838 249200 130844 249212
rect 6236 249172 130844 249200
rect 6236 249160 6242 249172
rect 130838 249160 130844 249172
rect 130896 249160 130902 249212
rect 191098 249160 191104 249212
rect 191156 249200 191162 249212
rect 359458 249200 359464 249212
rect 191156 249172 359464 249200
rect 191156 249160 191162 249172
rect 359458 249160 359464 249172
rect 359516 249160 359522 249212
rect 96982 249092 96988 249144
rect 97040 249132 97046 249144
rect 479518 249132 479524 249144
rect 97040 249104 479524 249132
rect 97040 249092 97046 249104
rect 479518 249092 479524 249104
rect 479576 249092 479582 249144
rect 85666 249024 85672 249076
rect 85724 249064 85730 249076
rect 545758 249064 545764 249076
rect 85724 249036 545764 249064
rect 85724 249024 85730 249036
rect 545758 249024 545764 249036
rect 545816 249024 545822 249076
rect 59262 247868 59268 247920
rect 59320 247908 59326 247920
rect 187326 247908 187332 247920
rect 59320 247880 187332 247908
rect 59320 247868 59326 247880
rect 187326 247868 187332 247880
rect 187384 247868 187390 247920
rect 62022 247800 62028 247852
rect 62080 247840 62086 247852
rect 241790 247840 241796 247852
rect 62080 247812 241796 247840
rect 62080 247800 62086 247812
rect 241790 247800 241796 247812
rect 241848 247800 241854 247852
rect 38102 247732 38108 247784
rect 38160 247772 38166 247784
rect 261478 247772 261484 247784
rect 38160 247744 261484 247772
rect 38160 247732 38166 247744
rect 261478 247732 261484 247744
rect 261536 247732 261542 247784
rect 31570 247664 31576 247716
rect 31628 247704 31634 247716
rect 358814 247704 358820 247716
rect 31628 247676 358820 247704
rect 31628 247664 31634 247676
rect 358814 247664 358820 247676
rect 358872 247664 358878 247716
rect 95694 246984 95700 247036
rect 95752 247024 95758 247036
rect 207658 247024 207664 247036
rect 95752 246996 207664 247024
rect 95752 246984 95758 246996
rect 207658 246984 207664 246996
rect 207716 246984 207722 247036
rect 88242 246916 88248 246968
rect 88300 246956 88306 246968
rect 204898 246956 204904 246968
rect 88300 246928 204904 246956
rect 88300 246916 88306 246928
rect 204898 246916 204904 246928
rect 204956 246916 204962 246968
rect 8202 246848 8208 246900
rect 8260 246888 8266 246900
rect 128354 246888 128360 246900
rect 8260 246860 128360 246888
rect 8260 246848 8266 246860
rect 128354 246848 128360 246860
rect 128412 246848 128418 246900
rect 139302 246848 139308 246900
rect 139360 246888 139366 246900
rect 240686 246888 240692 246900
rect 139360 246860 240692 246888
rect 139360 246848 139366 246860
rect 240686 246848 240692 246860
rect 240744 246848 240750 246900
rect 111702 246780 111708 246832
rect 111760 246820 111766 246832
rect 240594 246820 240600 246832
rect 111760 246792 240600 246820
rect 111760 246780 111766 246792
rect 240594 246780 240600 246792
rect 240652 246780 240658 246832
rect 36814 246712 36820 246764
rect 36872 246752 36878 246764
rect 107654 246752 107660 246764
rect 36872 246724 107660 246752
rect 36872 246712 36878 246724
rect 107654 246712 107660 246724
rect 107712 246712 107718 246764
rect 114554 246712 114560 246764
rect 114612 246752 114618 246764
rect 282914 246752 282920 246764
rect 114612 246724 282920 246752
rect 114612 246712 114618 246724
rect 282914 246712 282920 246724
rect 282972 246712 282978 246764
rect 3694 246644 3700 246696
rect 3752 246684 3758 246696
rect 152182 246684 152188 246696
rect 3752 246656 152188 246684
rect 3752 246644 3758 246656
rect 152182 246644 152188 246656
rect 152240 246644 152246 246696
rect 218146 246644 218152 246696
rect 218204 246684 218210 246696
rect 412634 246684 412640 246696
rect 218204 246656 412640 246684
rect 218204 246644 218210 246656
rect 412634 246644 412640 246656
rect 412692 246644 412698 246696
rect 34054 246576 34060 246628
rect 34112 246616 34118 246628
rect 372706 246616 372712 246628
rect 34112 246588 372712 246616
rect 34112 246576 34118 246588
rect 372706 246576 372712 246588
rect 372764 246576 372770 246628
rect 103238 246508 103244 246560
rect 103296 246548 103302 246560
rect 477494 246548 477500 246560
rect 103296 246520 477500 246548
rect 103296 246508 103302 246520
rect 477494 246508 477500 246520
rect 477552 246508 477558 246560
rect 76926 246440 76932 246492
rect 76984 246480 76990 246492
rect 486418 246480 486424 246492
rect 76984 246452 486424 246480
rect 76984 246440 76990 246452
rect 486418 246440 486424 246452
rect 486476 246440 486482 246492
rect 73154 246372 73160 246424
rect 73212 246412 73218 246424
rect 485038 246412 485044 246424
rect 73212 246384 485044 246412
rect 73212 246372 73218 246384
rect 485038 246372 485044 246384
rect 485096 246372 485102 246424
rect 35066 246304 35072 246356
rect 35124 246344 35130 246356
rect 70486 246344 70492 246356
rect 35124 246316 70492 246344
rect 35124 246304 35130 246316
rect 70486 246304 70492 246316
rect 70544 246304 70550 246356
rect 99466 246304 99472 246356
rect 99524 246344 99530 246356
rect 542354 246344 542360 246356
rect 99524 246316 542360 246344
rect 99524 246304 99530 246316
rect 542354 246304 542360 246316
rect 542412 246304 542418 246356
rect 33778 246236 33784 246288
rect 33836 246276 33842 246288
rect 143442 246276 143448 246288
rect 33836 246248 143448 246276
rect 33836 246236 33842 246248
rect 143442 246236 143448 246248
rect 143500 246236 143506 246288
rect 24762 246168 24768 246220
rect 24820 246208 24826 246220
rect 129642 246208 129648 246220
rect 24820 246180 129648 246208
rect 24820 246168 24826 246180
rect 129642 246168 129648 246180
rect 129700 246168 129706 246220
rect 118326 246100 118332 246152
rect 118384 246140 118390 246152
rect 218054 246140 218060 246152
rect 118384 246112 218060 246140
rect 118384 246100 118390 246112
rect 218054 246100 218060 246112
rect 218112 246100 218118 246152
rect 35158 245284 35164 245336
rect 35216 245324 35222 245336
rect 134610 245324 134616 245336
rect 35216 245296 134616 245324
rect 35216 245284 35222 245296
rect 134610 245284 134616 245296
rect 134668 245284 134674 245336
rect 31018 245216 31024 245268
rect 31076 245256 31082 245268
rect 138382 245256 138388 245268
rect 31076 245228 138388 245256
rect 31076 245216 31082 245228
rect 138382 245216 138388 245228
rect 138440 245216 138446 245268
rect 115842 245148 115848 245200
rect 115900 245188 115906 245200
rect 234614 245188 234620 245200
rect 115900 245160 234620 245188
rect 115900 245148 115906 245160
rect 234614 245148 234620 245160
rect 234672 245148 234678 245200
rect 13078 245080 13084 245132
rect 13136 245120 13142 245132
rect 145926 245120 145932 245132
rect 13136 245092 145932 245120
rect 13136 245080 13142 245092
rect 145926 245080 145932 245092
rect 145984 245080 145990 245132
rect 33778 245012 33784 245064
rect 33836 245052 33842 245064
rect 168466 245052 168472 245064
rect 33836 245024 168472 245052
rect 33836 245012 33842 245024
rect 168466 245012 168472 245024
rect 168524 245012 168530 245064
rect 112070 244944 112076 244996
rect 112128 244984 112134 244996
rect 299474 244984 299480 244996
rect 112128 244956 299480 244984
rect 112128 244944 112134 244956
rect 299474 244944 299480 244956
rect 299532 244944 299538 244996
rect 35250 244876 35256 244928
rect 35308 244916 35314 244928
rect 172238 244916 172244 244928
rect 35308 244888 172244 244916
rect 35308 244876 35314 244888
rect 172238 244876 172244 244888
rect 172296 244876 172302 244928
rect 223666 244876 223672 244928
rect 223724 244916 223730 244928
rect 420178 244916 420184 244928
rect 223724 244888 420184 244916
rect 223724 244876 223730 244888
rect 420178 244876 420184 244888
rect 420236 244876 420242 244928
rect 25498 244808 25504 244860
rect 25556 244848 25562 244860
rect 164694 244848 164700 244860
rect 25556 244820 164700 244848
rect 25556 244808 25562 244820
rect 164694 244808 164700 244820
rect 164752 244808 164758 244860
rect 28258 244740 28264 244792
rect 28316 244780 28322 244792
rect 176010 244780 176016 244792
rect 28316 244752 176016 244780
rect 28316 244740 28322 244752
rect 176010 244740 176016 244752
rect 176068 244740 176074 244792
rect 6178 244672 6184 244724
rect 6236 244712 6242 244724
rect 179782 244712 179788 244724
rect 6236 244684 179788 244712
rect 6236 244672 6242 244684
rect 179782 244672 179788 244684
rect 179840 244672 179846 244724
rect 59354 244604 59360 244656
rect 59412 244644 59418 244656
rect 265618 244644 265624 244656
rect 59412 244616 265624 244644
rect 59412 244604 59418 244616
rect 265618 244604 265624 244616
rect 265676 244604 265682 244656
rect 55582 244536 55588 244588
rect 55640 244576 55646 244588
rect 262858 244576 262864 244588
rect 55640 244548 262864 244576
rect 55640 244536 55646 244548
rect 262858 244536 262864 244548
rect 262916 244536 262922 244588
rect 51810 244468 51816 244520
rect 51868 244508 51874 244520
rect 261478 244508 261484 244520
rect 51868 244480 261484 244508
rect 51868 244468 51874 244480
rect 261478 244468 261484 244480
rect 261536 244468 261542 244520
rect 48038 244400 48044 244452
rect 48096 244440 48102 244452
rect 258718 244440 258724 244452
rect 48096 244412 258724 244440
rect 48096 244400 48102 244412
rect 258718 244400 258724 244412
rect 258776 244400 258782 244452
rect 44266 244332 44272 244384
rect 44324 244372 44330 244384
rect 255958 244372 255964 244384
rect 44324 244344 255964 244372
rect 44324 244332 44330 244344
rect 255958 244332 255964 244344
rect 256016 244332 256022 244384
rect 100754 244264 100760 244316
rect 100812 244304 100818 244316
rect 579798 244304 579804 244316
rect 100812 244276 579804 244304
rect 100812 244264 100818 244276
rect 579798 244264 579804 244276
rect 579856 244264 579862 244316
rect 68094 244196 68100 244248
rect 68152 244236 68158 244248
rect 68830 244236 68836 244248
rect 68152 244208 68836 244236
rect 68152 244196 68158 244208
rect 68830 244196 68836 244208
rect 68888 244196 68894 244248
rect 69382 244196 69388 244248
rect 69440 244236 69446 244248
rect 70302 244236 70308 244248
rect 69440 244208 70308 244236
rect 69440 244196 69446 244208
rect 70302 244196 70308 244208
rect 70360 244196 70366 244248
rect 70670 244196 70676 244248
rect 70728 244236 70734 244248
rect 71682 244236 71688 244248
rect 70728 244208 71688 244236
rect 70728 244196 70734 244208
rect 71682 244196 71688 244208
rect 71740 244196 71746 244248
rect 71866 244196 71872 244248
rect 71924 244236 71930 244248
rect 73062 244236 73068 244248
rect 71924 244208 73068 244236
rect 71924 244196 71930 244208
rect 73062 244196 73068 244208
rect 73120 244196 73126 244248
rect 84470 244196 84476 244248
rect 84528 244236 84534 244248
rect 85482 244236 85488 244248
rect 84528 244208 85488 244236
rect 84528 244196 84534 244208
rect 85482 244196 85488 244208
rect 85540 244196 85546 244248
rect 86954 244196 86960 244248
rect 87012 244236 87018 244248
rect 88150 244236 88156 244248
rect 87012 244208 88156 244236
rect 87012 244196 87018 244208
rect 88150 244196 88156 244208
rect 88208 244196 88214 244248
rect 98270 244196 98276 244248
rect 98328 244236 98334 244248
rect 100018 244236 100024 244248
rect 98328 244208 100024 244236
rect 98328 244196 98334 244208
rect 100018 244196 100024 244208
rect 100076 244196 100082 244248
rect 110782 244196 110788 244248
rect 110840 244236 110846 244248
rect 111610 244236 111616 244248
rect 110840 244208 111616 244236
rect 110840 244196 110846 244208
rect 111610 244196 111616 244208
rect 111668 244196 111674 244248
rect 113266 244196 113272 244248
rect 113324 244236 113330 244248
rect 114462 244236 114468 244248
rect 113324 244208 114468 244236
rect 113324 244196 113330 244208
rect 114462 244196 114468 244208
rect 114520 244196 114526 244248
rect 117038 244196 117044 244248
rect 117096 244236 117102 244248
rect 117958 244236 117964 244248
rect 117096 244208 117964 244236
rect 117096 244196 117102 244208
rect 117958 244196 117964 244208
rect 118016 244196 118022 244248
rect 173158 244196 173164 244248
rect 173216 244236 173222 244248
rect 173216 244208 202276 244236
rect 173216 244196 173222 244208
rect 7558 244128 7564 244180
rect 7616 244168 7622 244180
rect 171042 244168 171048 244180
rect 7616 244140 171048 244168
rect 7616 244128 7622 244140
rect 171042 244128 171048 244140
rect 171100 244128 171106 244180
rect 171778 244128 171784 244180
rect 171836 244168 171842 244180
rect 202141 244171 202199 244177
rect 202141 244168 202153 244171
rect 171836 244140 202153 244168
rect 171836 244128 171842 244140
rect 202141 244137 202153 244140
rect 202187 244137 202199 244171
rect 202248 244168 202276 244208
rect 202322 244196 202328 244248
rect 202380 244236 202386 244248
rect 203518 244236 203524 244248
rect 202380 244208 203524 244236
rect 202380 244196 202386 244208
rect 203518 244196 203524 244208
rect 203576 244196 203582 244248
rect 208670 244196 208676 244248
rect 208728 244236 208734 244248
rect 209682 244236 209688 244248
rect 208728 244208 209688 244236
rect 208728 244196 208734 244208
rect 209682 244196 209688 244208
rect 209740 244196 209746 244248
rect 233694 244196 233700 244248
rect 233752 244236 233758 244248
rect 234522 244236 234528 244248
rect 233752 244208 234528 244236
rect 233752 244196 233758 244208
rect 234522 244196 234528 244208
rect 234580 244196 234586 244248
rect 238754 244196 238760 244248
rect 238812 244236 238818 244248
rect 240042 244236 240048 244248
rect 238812 244208 240048 244236
rect 238812 244196 238818 244208
rect 240042 244196 240048 244208
rect 240100 244196 240106 244248
rect 206094 244168 206100 244180
rect 202248 244140 206100 244168
rect 202141 244131 202199 244137
rect 206094 244128 206100 244140
rect 206152 244128 206158 244180
rect 213178 244128 213184 244180
rect 213236 244168 213242 244180
rect 213236 244140 226932 244168
rect 213236 244128 213242 244140
rect 169018 244060 169024 244112
rect 169076 244100 169082 244112
rect 222470 244100 222476 244112
rect 169076 244072 222476 244100
rect 169076 244060 169082 244072
rect 222470 244060 222476 244072
rect 222528 244060 222534 244112
rect 226904 244100 226932 244140
rect 226978 244128 226984 244180
rect 227036 244168 227042 244180
rect 236270 244168 236276 244180
rect 227036 244140 236276 244168
rect 227036 244128 227042 244140
rect 236270 244128 236276 244140
rect 236328 244128 236334 244180
rect 237466 244128 237472 244180
rect 237524 244168 237530 244180
rect 373258 244168 373264 244180
rect 237524 244140 373264 244168
rect 237524 244128 237530 244140
rect 373258 244128 373264 244140
rect 373316 244128 373322 244180
rect 228726 244100 228732 244112
rect 226904 244072 228732 244100
rect 228726 244060 228732 244072
rect 228784 244060 228790 244112
rect 229922 244060 229928 244112
rect 229980 244100 229986 244112
rect 377398 244100 377404 244112
rect 229980 244072 377404 244100
rect 229980 244060 229986 244072
rect 377398 244060 377404 244072
rect 377456 244060 377462 244112
rect 162118 243992 162124 244044
rect 162176 244032 162182 244044
rect 219894 244032 219900 244044
rect 162176 244004 219900 244032
rect 162176 243992 162182 244004
rect 219894 243992 219900 244004
rect 219952 243992 219958 244044
rect 224954 243992 224960 244044
rect 225012 244032 225018 244044
rect 385678 244032 385684 244044
rect 225012 244004 385684 244032
rect 225012 243992 225018 244004
rect 385678 243992 385684 244004
rect 385736 243992 385742 244044
rect 153838 243924 153844 243976
rect 153896 243964 153902 243976
rect 153896 243936 180794 243964
rect 153896 243924 153902 243936
rect 123294 243856 123300 243908
rect 123352 243896 123358 243908
rect 176838 243896 176844 243908
rect 123352 243868 176844 243896
rect 123352 243856 123358 243868
rect 176838 243856 176844 243868
rect 176896 243856 176902 243908
rect 180766 243896 180794 243936
rect 192294 243924 192300 243976
rect 192352 243964 192358 243976
rect 193122 243964 193128 243976
rect 192352 243936 193128 243964
rect 192352 243924 192358 243936
rect 193122 243924 193128 243936
rect 193180 243924 193186 243976
rect 197354 243924 197360 243976
rect 197412 243964 197418 243976
rect 198642 243964 198648 243976
rect 197412 243936 198648 243964
rect 197412 243924 197418 243936
rect 198642 243924 198648 243936
rect 198700 243924 198706 243976
rect 200758 243924 200764 243976
rect 200816 243964 200822 243976
rect 213638 243964 213644 243976
rect 200816 243936 213644 243964
rect 200816 243924 200822 243936
rect 213638 243924 213644 243936
rect 213696 243924 213702 243976
rect 214926 243924 214932 243976
rect 214984 243964 214990 243976
rect 380894 243964 380900 243976
rect 214984 243936 380900 243964
rect 214984 243924 214990 243936
rect 380894 243924 380900 243936
rect 380952 243924 380958 243976
rect 196066 243896 196072 243908
rect 180766 243868 196072 243896
rect 196066 243856 196072 243868
rect 196124 243856 196130 243908
rect 202141 243899 202199 243905
rect 202141 243865 202153 243899
rect 202187 243896 202199 243899
rect 207382 243896 207388 243908
rect 202187 243868 207388 243896
rect 202187 243865 202199 243868
rect 202141 243859 202199 243865
rect 207382 243856 207388 243868
rect 207440 243856 207446 243908
rect 211154 243856 211160 243908
rect 211212 243896 211218 243908
rect 218977 243899 219035 243905
rect 211212 243868 218928 243896
rect 211212 243856 211218 243868
rect 122098 243788 122104 243840
rect 122156 243828 122162 243840
rect 176746 243828 176752 243840
rect 122156 243800 176752 243828
rect 122156 243788 122162 243800
rect 176746 243788 176752 243800
rect 176804 243788 176810 243840
rect 214558 243788 214564 243840
rect 214616 243828 214622 243840
rect 218698 243828 218704 243840
rect 214616 243800 218704 243828
rect 214616 243788 214622 243800
rect 218698 243788 218704 243800
rect 218756 243788 218762 243840
rect 63126 243720 63132 243772
rect 63184 243760 63190 243772
rect 100754 243760 100760 243772
rect 63184 243732 100760 243760
rect 63184 243720 63190 243732
rect 100754 243720 100760 243732
rect 100812 243720 100818 243772
rect 120810 243720 120816 243772
rect 120868 243760 120874 243772
rect 176654 243760 176660 243772
rect 120868 243732 176660 243760
rect 120868 243720 120874 243732
rect 176654 243720 176660 243732
rect 176712 243720 176718 243772
rect 177298 243720 177304 243772
rect 177356 243760 177362 243772
rect 194870 243760 194876 243772
rect 177356 243732 194876 243760
rect 177356 243720 177362 243732
rect 194870 243720 194876 243732
rect 194928 243720 194934 243772
rect 195238 243720 195244 243772
rect 195296 243760 195302 243772
rect 204898 243760 204904 243772
rect 195296 243732 204904 243760
rect 195296 243720 195302 243732
rect 204898 243720 204904 243732
rect 204956 243720 204962 243772
rect 218900 243760 218928 243868
rect 218977 243865 218989 243899
rect 219023 243896 219035 243899
rect 376846 243896 376852 243908
rect 219023 243868 376852 243896
rect 219023 243865 219035 243868
rect 218977 243859 219035 243865
rect 376846 243856 376852 243868
rect 376904 243856 376910 243908
rect 219069 243831 219127 243837
rect 219069 243797 219081 243831
rect 219115 243828 219127 243831
rect 379606 243828 379612 243840
rect 219115 243800 379612 243828
rect 219115 243797 219127 243800
rect 219069 243791 219127 243797
rect 379606 243788 379612 243800
rect 379664 243788 379670 243840
rect 379514 243760 379520 243772
rect 218900 243732 379520 243760
rect 379514 243720 379520 243732
rect 379572 243720 379578 243772
rect 39666 243652 39672 243704
rect 39724 243692 39730 243704
rect 124582 243692 124588 243704
rect 39724 243664 124588 243692
rect 39724 243652 39730 243664
rect 124582 243652 124588 243664
rect 124640 243652 124646 243704
rect 131758 243652 131764 243704
rect 131816 243692 131822 243704
rect 198642 243692 198648 243704
rect 131816 243664 198648 243692
rect 131816 243652 131822 243664
rect 198642 243652 198648 243664
rect 198700 243652 198706 243704
rect 203610 243652 203616 243704
rect 203668 243692 203674 243704
rect 373994 243692 374000 243704
rect 203668 243664 374000 243692
rect 203668 243652 203674 243664
rect 373994 243652 374000 243664
rect 374052 243652 374058 243704
rect 39850 243584 39856 243636
rect 39908 243624 39914 243636
rect 125870 243624 125876 243636
rect 39908 243596 125876 243624
rect 39908 243584 39914 243596
rect 125870 243584 125876 243596
rect 125928 243584 125934 243636
rect 188522 243584 188528 243636
rect 188580 243624 188586 243636
rect 363046 243624 363052 243636
rect 188580 243596 363052 243624
rect 188580 243584 188586 243596
rect 363046 243584 363052 243596
rect 363104 243584 363110 243636
rect 36630 243516 36636 243568
rect 36688 243556 36694 243568
rect 132586 243556 132592 243568
rect 36688 243528 132592 243556
rect 36688 243516 36694 243528
rect 132586 243516 132592 243528
rect 132644 243516 132650 243568
rect 186038 243516 186044 243568
rect 186096 243556 186102 243568
rect 362954 243556 362960 243568
rect 186096 243528 362960 243556
rect 186096 243516 186102 243528
rect 362954 243516 362960 243528
rect 363012 243516 363018 243568
rect 60642 243448 60648 243500
rect 60700 243488 60706 243500
rect 115934 243488 115940 243500
rect 60700 243460 115940 243488
rect 60700 243448 60706 243460
rect 115934 243448 115940 243460
rect 115992 243448 115998 243500
rect 167638 243448 167644 243500
rect 167696 243488 167702 243500
rect 201126 243488 201132 243500
rect 167696 243460 201132 243488
rect 167696 243448 167702 243460
rect 201126 243448 201132 243460
rect 201184 243448 201190 243500
rect 209866 243448 209872 243500
rect 209924 243488 209930 243500
rect 218977 243491 219035 243497
rect 218977 243488 218989 243491
rect 209924 243460 218989 243488
rect 209924 243448 209930 243460
rect 218977 243457 218989 243460
rect 219023 243457 219035 243491
rect 218977 243451 219035 243457
rect 225598 243448 225604 243500
rect 225656 243488 225662 243500
rect 232222 243488 232228 243500
rect 225656 243460 232228 243488
rect 225656 243448 225662 243460
rect 232222 243448 232228 243460
rect 232280 243448 232286 243500
rect 61838 243380 61844 243432
rect 61896 243420 61902 243432
rect 184658 243420 184664 243432
rect 61896 243392 184664 243420
rect 61896 243380 61902 243392
rect 184658 243380 184664 243392
rect 184716 243380 184722 243432
rect 199838 243380 199844 243432
rect 199896 243420 199902 243432
rect 229738 243420 229744 243432
rect 199896 243392 229744 243420
rect 199896 243380 199902 243392
rect 229738 243380 229744 243392
rect 229796 243380 229802 243432
rect 46842 243312 46848 243364
rect 46900 243352 46906 243364
rect 172422 243352 172428 243364
rect 46900 243324 172428 243352
rect 46900 243312 46906 243324
rect 172422 243312 172428 243324
rect 172480 243312 172486 243364
rect 183554 243312 183560 243364
rect 183612 243352 183618 243364
rect 184842 243352 184848 243364
rect 183612 243324 184848 243352
rect 183612 243312 183618 243324
rect 184842 243312 184848 243324
rect 184900 243312 184906 243364
rect 212442 243312 212448 243364
rect 212500 243352 212506 243364
rect 219069 243355 219127 243361
rect 219069 243352 219081 243355
rect 212500 243324 219081 243352
rect 212500 243312 212506 243324
rect 219069 243321 219081 243324
rect 219115 243321 219127 243355
rect 219069 243315 219127 243321
rect 222838 243312 222844 243364
rect 222896 243352 222902 243364
rect 226242 243352 226248 243364
rect 222896 243324 226248 243352
rect 222896 243312 222902 243324
rect 226242 243312 226248 243324
rect 226300 243312 226306 243364
rect 31754 243244 31760 243296
rect 31812 243284 31818 243296
rect 162210 243284 162216 243296
rect 31812 243256 162216 243284
rect 31812 243244 31818 243256
rect 162210 243244 162216 243256
rect 162268 243244 162274 243296
rect 58066 243176 58072 243228
rect 58124 243216 58130 243228
rect 187694 243216 187700 243228
rect 58124 243188 187700 243216
rect 58124 243176 58130 243188
rect 187694 243176 187700 243188
rect 187752 243176 187758 243228
rect 232498 243176 232504 243228
rect 232556 243216 232562 243228
rect 234982 243216 234988 243228
rect 232556 243188 234988 243216
rect 232556 243176 232562 243188
rect 234982 243176 234988 243188
rect 235040 243176 235046 243228
rect 19978 243108 19984 243160
rect 20036 243148 20042 243160
rect 167270 243148 167276 243160
rect 20036 243120 167276 243148
rect 20036 243108 20042 243120
rect 167270 243108 167276 243120
rect 167328 243108 167334 243160
rect 13078 243040 13084 243092
rect 13136 243080 13142 243092
rect 174722 243080 174728 243092
rect 13136 243052 174728 243080
rect 13136 243040 13142 243052
rect 174722 243040 174728 243052
rect 174780 243040 174786 243092
rect 220078 243040 220084 243092
rect 220136 243080 220142 243092
rect 227438 243080 227444 243092
rect 220136 243052 227444 243080
rect 220136 243040 220142 243052
rect 227438 243040 227444 243052
rect 227496 243040 227502 243092
rect 15838 242972 15844 243024
rect 15896 243012 15902 243024
rect 178494 243012 178500 243024
rect 15896 242984 178500 243012
rect 15896 242972 15902 242984
rect 178494 242972 178500 242984
rect 178552 242972 178558 243024
rect 36538 242904 36544 242956
rect 36596 242944 36602 242956
rect 40586 242944 40592 242956
rect 36596 242916 40592 242944
rect 36596 242904 36602 242916
rect 40586 242904 40592 242916
rect 40644 242904 40650 242956
rect 100754 242904 100760 242956
rect 100812 242944 100818 242956
rect 102042 242944 102048 242956
rect 100812 242916 102048 242944
rect 100812 242904 100818 242916
rect 102042 242904 102048 242916
rect 102100 242904 102106 242956
rect 38562 242836 38568 242888
rect 38620 242876 38626 242888
rect 39298 242876 39304 242888
rect 38620 242848 39304 242876
rect 38620 242836 38626 242848
rect 39298 242836 39304 242848
rect 39356 242836 39362 242888
rect 39850 242836 39856 242888
rect 39908 242876 39914 242888
rect 91186 242876 91192 242888
rect 39908 242848 91192 242876
rect 39908 242836 39914 242848
rect 91186 242836 91192 242848
rect 91244 242836 91250 242888
rect 92382 242836 92388 242888
rect 92440 242876 92446 242888
rect 240226 242876 240232 242888
rect 92440 242848 240232 242876
rect 92440 242836 92446 242848
rect 240226 242836 240232 242848
rect 240284 242836 240290 242888
rect 32766 242768 32772 242820
rect 32824 242808 32830 242820
rect 70578 242808 70584 242820
rect 32824 242780 70584 242808
rect 32824 242768 32830 242780
rect 70578 242768 70584 242780
rect 70636 242768 70642 242820
rect 82722 242768 82728 242820
rect 82780 242808 82786 242820
rect 243354 242808 243360 242820
rect 82780 242780 243360 242808
rect 82780 242768 82786 242780
rect 243354 242768 243360 242780
rect 243412 242768 243418 242820
rect 68922 242700 68928 242752
rect 68980 242740 68986 242752
rect 243262 242740 243268 242752
rect 68980 242712 243268 242740
rect 68980 242700 68986 242712
rect 243262 242700 243268 242712
rect 243320 242700 243326 242752
rect 63402 242632 63408 242684
rect 63460 242672 63466 242684
rect 240318 242672 240324 242684
rect 63460 242644 240324 242672
rect 63460 242632 63466 242644
rect 240318 242632 240324 242644
rect 240376 242632 240382 242684
rect 32950 242564 32956 242616
rect 33008 242604 33014 242616
rect 337562 242604 337568 242616
rect 33008 242576 337568 242604
rect 33008 242564 33014 242576
rect 337562 242564 337568 242576
rect 337620 242564 337626 242616
rect 35526 242496 35532 242548
rect 35584 242536 35590 242548
rect 376754 242536 376760 242548
rect 35584 242508 376760 242536
rect 35584 242496 35590 242508
rect 376754 242496 376760 242508
rect 376812 242496 376818 242548
rect 36446 242428 36452 242480
rect 36504 242468 36510 242480
rect 385034 242468 385040 242480
rect 36504 242440 385040 242468
rect 36504 242428 36510 242440
rect 385034 242428 385040 242440
rect 385092 242428 385098 242480
rect 35342 242360 35348 242412
rect 35400 242400 35406 242412
rect 420914 242400 420920 242412
rect 35400 242372 420920 242400
rect 35400 242360 35406 242372
rect 420914 242360 420920 242372
rect 420972 242360 420978 242412
rect 37182 242292 37188 242344
rect 37240 242332 37246 242344
rect 440234 242332 440240 242344
rect 37240 242304 440240 242332
rect 37240 242292 37246 242304
rect 440234 242292 440240 242304
rect 440292 242292 440298 242344
rect 39206 242224 39212 242276
rect 39264 242264 39270 242276
rect 442994 242264 443000 242276
rect 39264 242236 443000 242264
rect 39264 242224 39270 242236
rect 442994 242224 443000 242236
rect 443052 242224 443058 242276
rect 3418 242156 3424 242208
rect 3476 242196 3482 242208
rect 31754 242196 31760 242208
rect 3476 242168 31760 242196
rect 3476 242156 3482 242168
rect 31754 242156 31760 242168
rect 31812 242156 31818 242208
rect 64782 242156 64788 242208
rect 64840 242196 64846 242208
rect 244366 242196 244372 242208
rect 64840 242168 244372 242196
rect 64840 242156 64846 242168
rect 244366 242156 244372 242168
rect 244424 242156 244430 242208
rect 39022 242088 39028 242140
rect 39080 242128 39086 242140
rect 88426 242128 88432 242140
rect 39080 242100 88432 242128
rect 39080 242088 39086 242100
rect 88426 242088 88432 242100
rect 88484 242088 88490 242140
rect 96338 242088 96344 242140
rect 96396 242128 96402 242140
rect 244274 242128 244280 242140
rect 96396 242100 244280 242128
rect 96396 242088 96402 242100
rect 244274 242088 244280 242100
rect 244332 242088 244338 242140
rect 39942 242020 39948 242072
rect 40000 242060 40006 242072
rect 97994 242060 98000 242072
rect 40000 242032 98000 242060
rect 40000 242020 40006 242032
rect 97994 242020 98000 242032
rect 98052 242020 98058 242072
rect 35618 241952 35624 242004
rect 35676 241992 35682 242004
rect 82906 241992 82912 242004
rect 35676 241964 82912 241992
rect 35676 241952 35682 241964
rect 82906 241952 82912 241964
rect 82964 241952 82970 242004
rect 34146 241884 34152 241936
rect 34204 241924 34210 241936
rect 69106 241924 69112 241936
rect 34204 241896 69112 241924
rect 34204 241884 34210 241896
rect 69106 241884 69112 241896
rect 69164 241884 69170 241936
rect 39114 241476 39120 241528
rect 39172 241516 39178 241528
rect 39850 241516 39856 241528
rect 39172 241488 39856 241516
rect 39172 241476 39178 241488
rect 39850 241476 39856 241488
rect 39908 241476 39914 241528
rect 24118 241408 24124 241460
rect 24176 241448 24182 241460
rect 173158 241448 173164 241460
rect 24176 241420 173164 241448
rect 24176 241408 24182 241420
rect 173158 241408 173164 241420
rect 173216 241408 173222 241460
rect 37826 241340 37832 241392
rect 37884 241380 37890 241392
rect 43438 241380 43444 241392
rect 37884 241352 43444 241380
rect 37884 241340 37890 241352
rect 43438 241340 43444 241352
rect 43496 241340 43502 241392
rect 38286 241272 38292 241324
rect 38344 241312 38350 241324
rect 48958 241312 48964 241324
rect 38344 241284 48964 241312
rect 38344 241272 38350 241284
rect 48958 241272 48964 241284
rect 49016 241272 49022 241324
rect 38562 241204 38568 241256
rect 38620 241244 38626 241256
rect 42058 241244 42064 241256
rect 38620 241216 42064 241244
rect 38620 241204 38626 241216
rect 42058 241204 42064 241216
rect 42116 241204 42122 241256
rect 50338 241244 50344 241256
rect 42260 241216 50344 241244
rect 38838 241136 38844 241188
rect 38896 241176 38902 241188
rect 42153 241179 42211 241185
rect 42153 241176 42165 241179
rect 38896 241148 42165 241176
rect 38896 241136 38902 241148
rect 42153 241145 42165 241148
rect 42199 241145 42211 241179
rect 42153 241139 42211 241145
rect 37734 241068 37740 241120
rect 37792 241108 37798 241120
rect 42260 241108 42288 241216
rect 50338 241204 50344 241216
rect 50396 241204 50402 241256
rect 57146 241244 57152 241256
rect 57107 241216 57152 241244
rect 57146 241204 57152 241216
rect 57204 241204 57210 241256
rect 42337 241179 42395 241185
rect 42337 241145 42349 241179
rect 42383 241176 42395 241179
rect 45922 241176 45928 241188
rect 42383 241148 45554 241176
rect 45883 241148 45928 241176
rect 42383 241145 42395 241148
rect 42337 241139 42395 241145
rect 43346 241108 43352 241120
rect 37792 241080 42288 241108
rect 43307 241080 43352 241108
rect 37792 241068 37798 241080
rect 43346 241068 43352 241080
rect 43404 241068 43410 241120
rect 45526 241108 45554 241148
rect 45922 241136 45928 241148
rect 45980 241136 45986 241188
rect 49602 241176 49608 241188
rect 49563 241148 49608 241176
rect 49602 241136 49608 241148
rect 49660 241136 49666 241188
rect 50890 241176 50896 241188
rect 50851 241148 50896 241176
rect 50890 241136 50896 241148
rect 50948 241136 50954 241188
rect 53466 241176 53472 241188
rect 53427 241148 53472 241176
rect 53466 241136 53472 241148
rect 53524 241136 53530 241188
rect 54570 241176 54576 241188
rect 54531 241148 54576 241176
rect 54570 241136 54576 241148
rect 54628 241136 54634 241188
rect 54665 241179 54723 241185
rect 54665 241145 54677 241179
rect 54711 241176 54723 241179
rect 64966 241176 64972 241188
rect 54711 241148 64972 241176
rect 54711 241145 54723 241148
rect 54665 241139 54723 241145
rect 64966 241136 64972 241148
rect 65024 241136 65030 241188
rect 115934 241176 115940 241188
rect 115895 241148 115940 241176
rect 115934 241136 115940 241148
rect 115992 241136 115998 241188
rect 236638 241136 236644 241188
rect 236696 241176 236702 241188
rect 241606 241176 241612 241188
rect 236696 241148 241612 241176
rect 236696 241136 236702 241148
rect 241606 241136 241612 241148
rect 241664 241136 241670 241188
rect 66346 241108 66352 241120
rect 45526 241080 66352 241108
rect 66346 241068 66352 241080
rect 66404 241068 66410 241120
rect 82998 241108 83004 241120
rect 82959 241080 83004 241108
rect 82998 241068 83004 241080
rect 83056 241068 83062 241120
rect 88058 241068 88064 241120
rect 88116 241108 88122 241120
rect 241882 241108 241888 241120
rect 88116 241080 241888 241108
rect 88116 241068 88122 241080
rect 241882 241068 241888 241080
rect 241940 241068 241946 241120
rect 32398 241000 32404 241052
rect 32456 241040 32462 241052
rect 165614 241040 165620 241052
rect 32456 241012 165620 241040
rect 32456 241000 32462 241012
rect 165614 241000 165620 241012
rect 165672 241000 165678 241052
rect 221458 241000 221464 241052
rect 221516 241040 221522 241052
rect 241698 241040 241704 241052
rect 221516 241012 241704 241040
rect 221516 241000 221522 241012
rect 241698 241000 241704 241012
rect 241756 241000 241762 241052
rect 31018 240932 31024 240984
rect 31076 240972 31082 240984
rect 169570 240972 169576 240984
rect 31076 240944 169576 240972
rect 31076 240932 31082 240944
rect 169570 240932 169576 240944
rect 169628 240932 169634 240984
rect 172422 240932 172428 240984
rect 172480 240972 172486 240984
rect 172480 240944 177160 240972
rect 172480 240932 172486 240944
rect 21358 240864 21364 240916
rect 21416 240904 21422 240916
rect 177022 240904 177028 240916
rect 21416 240876 177028 240904
rect 21416 240864 21422 240876
rect 177022 240864 177028 240876
rect 177080 240864 177086 240916
rect 38746 240796 38752 240848
rect 38804 240836 38810 240848
rect 54665 240839 54723 240845
rect 54665 240836 54677 240839
rect 38804 240808 54677 240836
rect 38804 240796 38810 240808
rect 54665 240805 54677 240808
rect 54711 240805 54723 240839
rect 177132 240836 177160 240944
rect 187694 240932 187700 240984
rect 187752 240972 187758 240984
rect 580350 240972 580356 240984
rect 187752 240944 580356 240972
rect 187752 240932 187758 240944
rect 580350 240932 580356 240944
rect 580408 240932 580414 240984
rect 180886 240904 180892 240916
rect 180847 240876 180892 240904
rect 180886 240864 180892 240876
rect 180944 240864 180950 240916
rect 182082 240904 182088 240916
rect 182043 240876 182088 240904
rect 182082 240864 182088 240876
rect 182140 240864 182146 240916
rect 184658 240864 184664 240916
rect 184716 240904 184722 240916
rect 580442 240904 580448 240916
rect 184716 240876 580448 240904
rect 184716 240864 184722 240876
rect 580442 240864 580448 240876
rect 580500 240864 580506 240916
rect 580258 240836 580264 240848
rect 177132 240808 580264 240836
rect 54665 240799 54723 240805
rect 580258 240796 580264 240808
rect 580316 240796 580322 240848
rect 38930 240728 38936 240780
rect 38988 240768 38994 240780
rect 83001 240771 83059 240777
rect 83001 240768 83013 240771
rect 38988 240740 83013 240768
rect 38988 240728 38994 240740
rect 83001 240737 83013 240740
rect 83047 240737 83059 240771
rect 83001 240731 83059 240737
rect 115937 240771 115995 240777
rect 115937 240737 115949 240771
rect 115983 240768 115995 240771
rect 579798 240768 579804 240780
rect 115983 240740 579804 240768
rect 115983 240737 115995 240740
rect 115937 240731 115995 240737
rect 579798 240728 579804 240740
rect 579856 240728 579862 240780
rect 14458 240660 14464 240712
rect 14516 240700 14522 240712
rect 182085 240703 182143 240709
rect 182085 240700 182097 240703
rect 14516 240672 182097 240700
rect 14516 240660 14522 240672
rect 182085 240669 182097 240672
rect 182131 240669 182143 240703
rect 182085 240663 182143 240669
rect 10318 240592 10324 240644
rect 10376 240632 10382 240644
rect 180889 240635 180947 240641
rect 180889 240632 180901 240635
rect 10376 240604 180901 240632
rect 10376 240592 10382 240604
rect 180889 240601 180901 240604
rect 180935 240601 180947 240635
rect 180889 240595 180947 240601
rect 57149 240567 57207 240573
rect 57149 240533 57161 240567
rect 57195 240564 57207 240567
rect 273898 240564 273904 240576
rect 57195 240536 273904 240564
rect 57195 240533 57207 240536
rect 57149 240527 57207 240533
rect 273898 240524 273904 240536
rect 273956 240524 273962 240576
rect 53469 240499 53527 240505
rect 53469 240465 53481 240499
rect 53515 240496 53527 240499
rect 272518 240496 272524 240508
rect 53515 240468 272524 240496
rect 53515 240465 53527 240468
rect 53469 240459 53527 240465
rect 272518 240456 272524 240468
rect 272576 240456 272582 240508
rect 49605 240431 49663 240437
rect 49605 240397 49617 240431
rect 49651 240428 49663 240431
rect 269758 240428 269764 240440
rect 49651 240400 269764 240428
rect 49651 240397 49663 240400
rect 49605 240391 49663 240397
rect 269758 240388 269764 240400
rect 269816 240388 269822 240440
rect 45925 240363 45983 240369
rect 45925 240329 45937 240363
rect 45971 240360 45983 240363
rect 268378 240360 268384 240372
rect 45971 240332 268384 240360
rect 45971 240329 45983 240332
rect 45925 240323 45983 240329
rect 268378 240320 268384 240332
rect 268436 240320 268442 240372
rect 54573 240295 54631 240301
rect 54573 240261 54585 240295
rect 54619 240292 54631 240295
rect 280798 240292 280804 240304
rect 54619 240264 280804 240292
rect 54619 240261 54631 240264
rect 54573 240255 54631 240261
rect 280798 240252 280804 240264
rect 280856 240252 280862 240304
rect 50893 240227 50951 240233
rect 50893 240193 50905 240227
rect 50939 240224 50951 240227
rect 279418 240224 279424 240236
rect 50939 240196 279424 240224
rect 50939 240193 50951 240196
rect 50893 240187 50951 240193
rect 279418 240184 279424 240196
rect 279476 240184 279482 240236
rect 43349 240159 43407 240165
rect 43349 240125 43361 240159
rect 43395 240156 43407 240159
rect 276658 240156 276664 240168
rect 43395 240128 276664 240156
rect 43395 240125 43407 240128
rect 43349 240119 43407 240125
rect 276658 240116 276664 240128
rect 276716 240116 276722 240168
rect 242802 234540 242808 234592
rect 242860 234580 242866 234592
rect 391290 234580 391296 234592
rect 242860 234552 391296 234580
rect 242860 234540 242866 234552
rect 391290 234540 391296 234552
rect 391348 234540 391354 234592
rect 242802 223524 242808 223576
rect 242860 223564 242866 223576
rect 367738 223564 367744 223576
rect 242860 223536 367744 223564
rect 242860 223524 242866 223536
rect 367738 223524 367744 223536
rect 367796 223524 367802 223576
rect 35802 217948 35808 218000
rect 35860 217988 35866 218000
rect 38010 217988 38016 218000
rect 35860 217960 38016 217988
rect 35860 217948 35866 217960
rect 38010 217948 38016 217960
rect 38068 217948 38074 218000
rect 242802 217948 242808 218000
rect 242860 217988 242866 218000
rect 388438 217988 388444 218000
rect 242860 217960 388444 217988
rect 242860 217948 242866 217960
rect 388438 217948 388444 217960
rect 388496 217948 388502 218000
rect 3326 215228 3332 215280
rect 3384 215268 3390 215280
rect 25498 215268 25504 215280
rect 3384 215240 25504 215268
rect 3384 215228 3390 215240
rect 25498 215228 25504 215240
rect 25556 215228 25562 215280
rect 241974 212372 241980 212424
rect 242032 212412 242038 212424
rect 243446 212412 243452 212424
rect 242032 212384 243452 212412
rect 242032 212372 242038 212384
rect 243446 212372 243452 212384
rect 243504 212372 243510 212424
rect 242526 208292 242532 208344
rect 242584 208332 242590 208344
rect 427814 208332 427820 208344
rect 242584 208304 427820 208332
rect 242584 208292 242590 208304
rect 427814 208292 427820 208304
rect 427872 208292 427878 208344
rect 265618 206932 265624 206984
rect 265676 206972 265682 206984
rect 579890 206972 579896 206984
rect 265676 206944 579896 206972
rect 265676 206932 265682 206944
rect 579890 206932 579896 206944
rect 579948 206932 579954 206984
rect 3418 202784 3424 202836
rect 3476 202824 3482 202836
rect 19978 202824 19984 202836
rect 3476 202796 19984 202824
rect 3476 202784 3482 202796
rect 19978 202784 19984 202796
rect 20036 202784 20042 202836
rect 242434 202784 242440 202836
rect 242492 202824 242498 202836
rect 387058 202824 387064 202836
rect 242492 202796 387064 202824
rect 242492 202784 242498 202796
rect 387058 202784 387064 202796
rect 387116 202784 387122 202836
rect 242342 197276 242348 197328
rect 242400 197316 242406 197328
rect 424318 197316 424324 197328
rect 242400 197288 424324 197316
rect 242400 197276 242406 197288
rect 424318 197276 424324 197288
rect 424376 197276 424382 197328
rect 35342 195916 35348 195968
rect 35400 195956 35406 195968
rect 38010 195956 38016 195968
rect 35400 195928 38016 195956
rect 35400 195916 35406 195928
rect 38010 195916 38016 195928
rect 38068 195916 38074 195968
rect 273898 193128 273904 193180
rect 273956 193168 273962 193180
rect 580166 193168 580172 193180
rect 273956 193140 580172 193168
rect 273956 193128 273962 193140
rect 580166 193128 580172 193140
rect 580224 193128 580230 193180
rect 31386 191768 31392 191820
rect 31444 191808 31450 191820
rect 38010 191808 38016 191820
rect 31444 191780 38016 191808
rect 31444 191768 31450 191780
rect 38010 191768 38016 191780
rect 38068 191768 38074 191820
rect 3418 188980 3424 189032
rect 3476 189020 3482 189032
rect 32398 189020 32404 189032
rect 3476 188992 32404 189020
rect 3476 188980 3482 188992
rect 32398 188980 32404 188992
rect 32456 188980 32462 189032
rect 36446 187620 36452 187672
rect 36504 187660 36510 187672
rect 37366 187660 37372 187672
rect 36504 187632 37372 187660
rect 36504 187620 36510 187632
rect 37366 187620 37372 187632
rect 37424 187620 37430 187672
rect 37826 186396 37832 186448
rect 37884 186436 37890 186448
rect 40494 186436 40500 186448
rect 37884 186408 40500 186436
rect 37884 186396 37890 186408
rect 40494 186396 40500 186408
rect 40552 186396 40558 186448
rect 37090 186328 37096 186380
rect 37148 186368 37154 186380
rect 37918 186368 37924 186380
rect 37148 186340 37924 186368
rect 37148 186328 37154 186340
rect 37918 186328 37924 186340
rect 37976 186328 37982 186380
rect 242802 186260 242808 186312
rect 242860 186300 242866 186312
rect 386414 186300 386420 186312
rect 242860 186272 386420 186300
rect 242860 186260 242866 186272
rect 386414 186260 386420 186272
rect 386472 186260 386478 186312
rect 38378 183472 38384 183524
rect 38436 183512 38442 183524
rect 39482 183512 39488 183524
rect 38436 183484 39488 183512
rect 38436 183472 38442 183484
rect 39482 183472 39488 183484
rect 39540 183472 39546 183524
rect 242802 180752 242808 180804
rect 242860 180792 242866 180804
rect 417418 180792 417424 180804
rect 242860 180764 417424 180792
rect 242860 180752 242866 180764
rect 417418 180752 417424 180764
rect 417476 180752 417482 180804
rect 32674 177964 32680 178016
rect 32732 178004 32738 178016
rect 38010 178004 38016 178016
rect 32732 177976 38016 178004
rect 32732 177964 32738 177976
rect 38010 177964 38016 177976
rect 38068 177964 38074 178016
rect 242802 175176 242808 175228
rect 242860 175216 242866 175228
rect 415394 175216 415400 175228
rect 242860 175188 415400 175216
rect 242860 175176 242866 175188
rect 415394 175176 415400 175188
rect 415452 175176 415458 175228
rect 35434 173340 35440 173392
rect 35492 173380 35498 173392
rect 38010 173380 38016 173392
rect 35492 173352 38016 173380
rect 35492 173340 35498 173352
rect 38010 173340 38016 173352
rect 38068 173340 38074 173392
rect 241882 169940 241888 169992
rect 241940 169980 241946 169992
rect 244458 169980 244464 169992
rect 241940 169952 244464 169980
rect 241940 169940 241946 169952
rect 244458 169940 244464 169952
rect 244516 169940 244522 169992
rect 33962 169668 33968 169720
rect 34020 169708 34026 169720
rect 38010 169708 38016 169720
rect 34020 169680 38016 169708
rect 34020 169668 34026 169680
rect 38010 169668 38016 169680
rect 38068 169668 38074 169720
rect 262858 166948 262864 167000
rect 262916 166988 262922 167000
rect 580166 166988 580172 167000
rect 262916 166960 580172 166988
rect 262916 166948 262922 166960
rect 580166 166948 580172 166960
rect 580224 166948 580230 167000
rect 3234 164160 3240 164212
rect 3292 164200 3298 164212
rect 33778 164200 33784 164212
rect 3292 164172 33784 164200
rect 3292 164160 3298 164172
rect 33778 164160 33784 164172
rect 33836 164160 33842 164212
rect 34330 161372 34336 161424
rect 34388 161412 34394 161424
rect 38010 161412 38016 161424
rect 34388 161384 38016 161412
rect 34388 161372 34394 161384
rect 38010 161372 38016 161384
rect 38068 161372 38074 161424
rect 241882 159400 241888 159452
rect 241940 159440 241946 159452
rect 243354 159440 243360 159452
rect 241940 159412 243360 159440
rect 241940 159400 241946 159412
rect 243354 159400 243360 159412
rect 243412 159400 243418 159452
rect 272518 153144 272524 153196
rect 272576 153184 272582 153196
rect 579798 153184 579804 153196
rect 272576 153156 579804 153184
rect 272576 153144 272582 153156
rect 579798 153144 579804 153156
rect 579856 153144 579862 153196
rect 35526 151716 35532 151768
rect 35584 151756 35590 151768
rect 38010 151756 38016 151768
rect 35584 151728 38016 151756
rect 35584 151716 35590 151728
rect 38010 151716 38016 151728
rect 38068 151716 38074 151768
rect 3418 150220 3424 150272
rect 3476 150260 3482 150272
rect 7558 150260 7564 150272
rect 3476 150232 7564 150260
rect 3476 150220 3482 150232
rect 7558 150220 7564 150232
rect 7616 150220 7622 150272
rect 242802 148996 242808 149048
rect 242860 149036 242866 149048
rect 405734 149036 405740 149048
rect 242860 149008 405740 149036
rect 242860 148996 242866 149008
rect 405734 148996 405740 149008
rect 405792 148996 405798 149048
rect 35710 147568 35716 147620
rect 35768 147608 35774 147620
rect 38010 147608 38016 147620
rect 35768 147580 38016 147608
rect 35768 147568 35774 147580
rect 38010 147568 38016 147580
rect 38068 147568 38074 147620
rect 241882 143420 241888 143472
rect 241940 143460 241946 143472
rect 244642 143460 244648 143472
rect 241940 143432 244648 143460
rect 241940 143420 241946 143432
rect 244642 143420 244648 143432
rect 244700 143420 244706 143472
rect 34054 139340 34060 139392
rect 34112 139380 34118 139392
rect 38010 139380 38016 139392
rect 34112 139352 38016 139380
rect 34112 139340 34118 139352
rect 38010 139340 38016 139352
rect 38068 139340 38074 139392
rect 280798 139340 280804 139392
rect 280856 139380 280862 139392
rect 580166 139380 580172 139392
rect 280856 139352 580172 139380
rect 280856 139340 280862 139352
rect 580166 139340 580172 139352
rect 580224 139340 580230 139392
rect 3234 137912 3240 137964
rect 3292 137952 3298 137964
rect 31018 137952 31024 137964
rect 3292 137924 31024 137952
rect 3292 137912 3298 137924
rect 31018 137912 31024 137924
rect 31076 137912 31082 137964
rect 32858 131044 32864 131096
rect 32916 131084 32922 131096
rect 38010 131084 38016 131096
rect 32916 131056 38016 131084
rect 32916 131044 32922 131056
rect 38010 131044 38016 131056
rect 38068 131044 38074 131096
rect 242250 128256 242256 128308
rect 242308 128296 242314 128308
rect 393406 128296 393412 128308
rect 242308 128268 393412 128296
rect 242308 128256 242314 128268
rect 393406 128256 393412 128268
rect 393464 128256 393470 128308
rect 261478 126896 261484 126948
rect 261536 126936 261542 126948
rect 580166 126936 580172 126948
rect 261536 126908 580172 126936
rect 261536 126896 261542 126908
rect 580166 126896 580172 126908
rect 580224 126896 580230 126948
rect 32766 125128 32772 125180
rect 32824 125168 32830 125180
rect 38010 125168 38016 125180
rect 32824 125140 38016 125168
rect 32824 125128 32830 125140
rect 38010 125128 38016 125140
rect 38068 125128 38074 125180
rect 241974 122544 241980 122596
rect 242032 122584 242038 122596
rect 245654 122584 245660 122596
rect 242032 122556 245660 122584
rect 242032 122544 242038 122556
rect 245654 122544 245660 122556
rect 245712 122544 245718 122596
rect 34146 121388 34152 121440
rect 34204 121428 34210 121440
rect 37918 121428 37924 121440
rect 34204 121400 37924 121428
rect 34204 121388 34210 121400
rect 37918 121388 37924 121400
rect 37976 121388 37982 121440
rect 38194 117920 38200 117972
rect 38252 117960 38258 117972
rect 39390 117960 39396 117972
rect 38252 117932 39396 117960
rect 38252 117920 38258 117932
rect 39390 117920 39396 117932
rect 39448 117920 39454 117972
rect 242802 117240 242808 117292
rect 242860 117280 242866 117292
rect 254578 117280 254584 117292
rect 242860 117252 254584 117280
rect 242860 117240 242866 117252
rect 254578 117240 254584 117252
rect 254636 117240 254642 117292
rect 35618 113092 35624 113144
rect 35676 113132 35682 113144
rect 38010 113132 38016 113144
rect 35676 113104 38016 113132
rect 35676 113092 35682 113104
rect 38010 113092 38016 113104
rect 38068 113092 38074 113144
rect 269758 113092 269764 113144
rect 269816 113132 269822 113144
rect 580166 113132 580172 113144
rect 269816 113104 580172 113132
rect 269816 113092 269822 113104
rect 580166 113092 580172 113104
rect 580224 113092 580230 113144
rect 3418 111732 3424 111784
rect 3476 111772 3482 111784
rect 35250 111772 35256 111784
rect 3476 111744 35256 111772
rect 3476 111732 3482 111744
rect 35250 111732 35256 111744
rect 35308 111732 35314 111784
rect 241882 111596 241888 111648
rect 241940 111636 241946 111648
rect 243262 111636 243268 111648
rect 241940 111608 243268 111636
rect 241940 111596 241946 111608
rect 243262 111596 243268 111608
rect 243320 111596 243326 111648
rect 34422 108944 34428 108996
rect 34480 108984 34486 108996
rect 37642 108984 37648 108996
rect 34480 108956 37648 108984
rect 34480 108944 34486 108956
rect 37642 108944 37648 108956
rect 37700 108944 37706 108996
rect 241882 107516 241888 107568
rect 241940 107556 241946 107568
rect 244550 107556 244556 107568
rect 241940 107528 244556 107556
rect 241940 107516 241946 107528
rect 244550 107516 244556 107528
rect 244608 107516 244614 107568
rect 279418 100648 279424 100700
rect 279476 100688 279482 100700
rect 580166 100688 580172 100700
rect 279476 100660 580172 100688
rect 279476 100648 279482 100660
rect 580166 100648 580172 100660
rect 580224 100648 580230 100700
rect 3418 97928 3424 97980
rect 3476 97968 3482 97980
rect 13078 97968 13084 97980
rect 3476 97940 13084 97968
rect 3476 97928 3482 97940
rect 13078 97928 13084 97940
rect 13136 97928 13142 97980
rect 242802 95956 242808 96008
rect 242860 95996 242866 96008
rect 250438 95996 250444 96008
rect 242860 95968 250444 95996
rect 242860 95956 242866 95968
rect 250438 95956 250444 95968
rect 250496 95956 250502 96008
rect 34238 95140 34244 95192
rect 34296 95180 34302 95192
rect 38010 95180 38016 95192
rect 34296 95152 38016 95180
rect 34296 95140 34302 95152
rect 38010 95140 38016 95152
rect 38068 95140 38074 95192
rect 31478 90992 31484 91044
rect 31536 91032 31542 91044
rect 38010 91032 38016 91044
rect 31536 91004 38016 91032
rect 31536 90992 31542 91004
rect 38010 90992 38016 91004
rect 38068 90992 38074 91044
rect 258718 86912 258724 86964
rect 258776 86952 258782 86964
rect 580166 86952 580172 86964
rect 258776 86924 580172 86952
rect 258776 86912 258782 86924
rect 580166 86912 580172 86924
rect 580224 86912 580230 86964
rect 3142 85484 3148 85536
rect 3200 85524 3206 85536
rect 24118 85524 24124 85536
rect 3200 85496 24124 85524
rect 3200 85484 3206 85496
rect 24118 85484 24124 85496
rect 24176 85484 24182 85536
rect 242250 79976 242256 80028
rect 242308 80016 242314 80028
rect 249058 80016 249064 80028
rect 242308 79988 249064 80016
rect 242308 79976 242314 79988
rect 249058 79976 249064 79988
rect 249116 79976 249122 80028
rect 30282 76916 30288 76968
rect 30340 76956 30346 76968
rect 38010 76956 38016 76968
rect 30340 76928 38016 76956
rect 30340 76916 30346 76928
rect 38010 76916 38016 76928
rect 38068 76916 38074 76968
rect 241514 74468 241520 74520
rect 241572 74508 241578 74520
rect 243170 74508 243176 74520
rect 241572 74480 243176 74508
rect 241572 74468 241578 74480
rect 243170 74468 243176 74480
rect 243228 74468 243234 74520
rect 268378 73108 268384 73160
rect 268436 73148 268442 73160
rect 579982 73148 579988 73160
rect 268436 73120 579988 73148
rect 268436 73108 268442 73120
rect 579982 73108 579988 73120
rect 580040 73108 580046 73160
rect 3418 71680 3424 71732
rect 3476 71720 3482 71732
rect 28258 71720 28264 71732
rect 3476 71692 28264 71720
rect 3476 71680 3482 71692
rect 28258 71680 28264 71692
rect 28316 71680 28322 71732
rect 31662 68960 31668 69012
rect 31720 69000 31726 69012
rect 38010 69000 38016 69012
rect 31720 68972 38016 69000
rect 31720 68960 31726 68972
rect 38010 68960 38016 68972
rect 38068 68960 38074 69012
rect 242802 64812 242808 64864
rect 242860 64852 242866 64864
rect 356146 64852 356152 64864
rect 242860 64824 356152 64852
rect 242860 64812 242866 64824
rect 356146 64812 356152 64824
rect 356204 64812 356210 64864
rect 31570 60664 31576 60716
rect 31628 60704 31634 60716
rect 38010 60704 38016 60716
rect 31628 60676 38016 60704
rect 31628 60664 31634 60676
rect 38010 60664 38016 60676
rect 38068 60664 38074 60716
rect 3050 59304 3056 59356
rect 3108 59344 3114 59356
rect 15838 59344 15844 59356
rect 3108 59316 15844 59344
rect 3108 59304 3114 59316
rect 15838 59304 15844 59316
rect 15896 59304 15902 59356
rect 241514 58896 241520 58948
rect 241572 58936 241578 58948
rect 244366 58936 244372 58948
rect 241572 58908 244372 58936
rect 241572 58896 241578 58908
rect 244366 58896 244372 58908
rect 244424 58896 244430 58948
rect 35066 56516 35072 56568
rect 35124 56556 35130 56568
rect 38010 56556 38016 56568
rect 35124 56528 38016 56556
rect 35124 56516 35130 56528
rect 38010 56516 38016 56528
rect 38068 56516 38074 56568
rect 241974 53728 241980 53780
rect 242032 53768 242038 53780
rect 357434 53768 357440 53780
rect 242032 53740 357440 53768
rect 242032 53728 242038 53740
rect 357434 53728 357440 53740
rect 357492 53728 357498 53780
rect 32950 46860 32956 46912
rect 33008 46900 33014 46912
rect 38010 46900 38016 46912
rect 33008 46872 38016 46900
rect 33008 46860 33014 46872
rect 38010 46860 38016 46872
rect 38068 46860 38074 46912
rect 255958 46860 255964 46912
rect 256016 46900 256022 46912
rect 580166 46900 580172 46912
rect 256016 46872 580172 46900
rect 256016 46860 256022 46872
rect 580166 46860 580172 46872
rect 580224 46860 580230 46912
rect 3418 45500 3424 45552
rect 3476 45540 3482 45552
rect 21358 45540 21364 45552
rect 3476 45512 21364 45540
rect 3476 45500 3482 45512
rect 21358 45500 21364 45512
rect 21416 45500 21422 45552
rect 33042 42712 33048 42764
rect 33100 42752 33106 42764
rect 38010 42752 38016 42764
rect 33100 42724 38016 42752
rect 33100 42712 33106 42724
rect 38010 42712 38016 42724
rect 38068 42712 38074 42764
rect 36538 39312 36544 39364
rect 36596 39352 36602 39364
rect 580258 39352 580264 39364
rect 36596 39324 580264 39352
rect 36596 39312 36602 39324
rect 580258 39312 580264 39324
rect 580316 39312 580322 39364
rect 220170 39040 220176 39092
rect 220228 39080 220234 39092
rect 355318 39080 355324 39092
rect 220228 39052 355324 39080
rect 220228 39040 220234 39052
rect 355318 39040 355324 39052
rect 355376 39040 355382 39092
rect 232958 38972 232964 39024
rect 233016 39012 233022 39024
rect 392578 39012 392584 39024
rect 233016 38984 392584 39012
rect 233016 38972 233022 38984
rect 392578 38972 392584 38984
rect 392636 38972 392642 39024
rect 200206 38904 200212 38956
rect 200264 38944 200270 38956
rect 367094 38944 367100 38956
rect 200264 38916 367100 38944
rect 200264 38904 200270 38916
rect 367094 38904 367100 38916
rect 367152 38904 367158 38956
rect 223022 38836 223028 38888
rect 223080 38876 223086 38888
rect 397546 38876 397552 38888
rect 223080 38848 397552 38876
rect 223080 38836 223086 38848
rect 397546 38836 397552 38848
rect 397604 38836 397610 38888
rect 225874 38768 225880 38820
rect 225932 38808 225938 38820
rect 402974 38808 402980 38820
rect 225932 38780 402980 38808
rect 225932 38768 225938 38780
rect 402974 38768 402980 38780
rect 403032 38768 403038 38820
rect 230106 38700 230112 38752
rect 230164 38740 230170 38752
rect 430574 38740 430580 38752
rect 230164 38712 430580 38740
rect 230164 38700 230170 38712
rect 430574 38700 430580 38712
rect 430632 38700 430638 38752
rect 38470 38632 38476 38684
rect 38528 38672 38534 38684
rect 215846 38672 215852 38684
rect 38528 38644 215852 38672
rect 38528 38632 38534 38644
rect 215846 38632 215852 38644
rect 215904 38632 215910 38684
rect 231578 38632 231584 38684
rect 231636 38672 231642 38684
rect 433334 38672 433340 38684
rect 231636 38644 433340 38672
rect 231636 38632 231642 38644
rect 433334 38632 433340 38644
rect 433392 38632 433398 38684
rect 39298 38564 39304 38616
rect 39356 38604 39362 38616
rect 40678 38604 40684 38616
rect 39356 38576 40684 38604
rect 39356 38564 39362 38576
rect 40678 38564 40684 38576
rect 40736 38604 40742 38616
rect 195882 38604 195888 38616
rect 40736 38576 195888 38604
rect 40736 38564 40742 38576
rect 195882 38564 195888 38576
rect 195940 38564 195946 38616
rect 237282 38564 237288 38616
rect 237340 38604 237346 38616
rect 244274 38604 244280 38616
rect 237340 38576 244280 38604
rect 237340 38564 237346 38576
rect 244274 38564 244280 38576
rect 244332 38564 244338 38616
rect 37090 38496 37096 38548
rect 37148 38536 37154 38548
rect 212994 38536 213000 38548
rect 37148 38508 213000 38536
rect 37148 38496 37154 38508
rect 212994 38496 213000 38508
rect 213052 38496 213058 38548
rect 224402 38496 224408 38548
rect 224460 38536 224466 38548
rect 239582 38536 239588 38548
rect 224460 38508 239588 38536
rect 224460 38496 224466 38508
rect 239582 38496 239588 38508
rect 239640 38496 239646 38548
rect 40402 38428 40408 38480
rect 40460 38468 40466 38480
rect 204438 38468 204444 38480
rect 40460 38440 204444 38468
rect 40460 38428 40466 38440
rect 204438 38428 204444 38440
rect 204496 38428 204502 38480
rect 227254 38428 227260 38480
rect 227312 38468 227318 38480
rect 240134 38468 240140 38480
rect 227312 38440 240140 38468
rect 227312 38428 227318 38440
rect 240134 38428 240140 38440
rect 240192 38428 240198 38480
rect 39482 38360 39488 38412
rect 39540 38400 39546 38412
rect 197354 38400 197360 38412
rect 39540 38372 197360 38400
rect 39540 38360 39546 38372
rect 197354 38360 197360 38372
rect 197412 38360 197418 38412
rect 228726 38360 228732 38412
rect 228784 38400 228790 38412
rect 240226 38400 240232 38412
rect 228784 38372 240232 38400
rect 228784 38360 228790 38372
rect 240226 38360 240232 38372
rect 240284 38360 240290 38412
rect 207290 38292 207296 38344
rect 207348 38332 207354 38344
rect 365714 38332 365720 38344
rect 207348 38304 365720 38332
rect 207348 38292 207354 38304
rect 365714 38292 365720 38304
rect 365772 38292 365778 38344
rect 59998 38224 60004 38276
rect 60056 38264 60062 38276
rect 69106 38264 69112 38276
rect 60056 38236 69112 38264
rect 60056 38224 60062 38236
rect 69106 38224 69112 38236
rect 69164 38224 69170 38276
rect 90358 38224 90364 38276
rect 90416 38264 90422 38276
rect 147490 38264 147496 38276
rect 90416 38236 147496 38264
rect 90416 38224 90422 38236
rect 147490 38224 147496 38236
rect 147548 38224 147554 38276
rect 151078 38224 151084 38276
rect 151136 38264 151142 38276
rect 160278 38264 160284 38276
rect 151136 38236 160284 38264
rect 151136 38224 151142 38236
rect 160278 38224 160284 38236
rect 160336 38224 160342 38276
rect 234430 38224 234436 38276
rect 234488 38264 234494 38276
rect 391198 38264 391204 38276
rect 234488 38236 391204 38264
rect 234488 38224 234494 38236
rect 391198 38224 391204 38236
rect 391256 38224 391262 38276
rect 66898 38156 66904 38208
rect 66956 38196 66962 38208
rect 79134 38196 79140 38208
rect 66956 38168 79140 38196
rect 66956 38156 66962 38168
rect 79134 38156 79140 38168
rect 79192 38156 79198 38208
rect 156046 38196 156052 38208
rect 103486 38168 156052 38196
rect 61378 38088 61384 38140
rect 61436 38128 61442 38140
rect 74810 38128 74816 38140
rect 61436 38100 74816 38128
rect 61436 38088 61442 38100
rect 74810 38088 74816 38100
rect 74868 38088 74874 38140
rect 79318 38088 79324 38140
rect 79376 38128 79382 38140
rect 91922 38128 91928 38140
rect 79376 38100 91928 38128
rect 79376 38088 79382 38100
rect 91922 38088 91928 38100
rect 91980 38088 91986 38140
rect 37090 38020 37096 38072
rect 37148 38060 37154 38072
rect 83366 38060 83372 38072
rect 37148 38032 83372 38060
rect 37148 38020 37154 38032
rect 83366 38020 83372 38032
rect 83424 38020 83430 38072
rect 39942 37952 39948 38004
rect 40000 37992 40006 38004
rect 87690 37992 87696 38004
rect 40000 37964 87696 37992
rect 40000 37952 40006 37964
rect 87690 37952 87696 37964
rect 87748 37952 87754 38004
rect 46842 37884 46848 37936
rect 46900 37924 46906 37936
rect 96154 37924 96160 37936
rect 46900 37896 96160 37924
rect 46900 37884 46906 37896
rect 96154 37884 96160 37896
rect 96212 37884 96218 37936
rect 100018 37884 100024 37936
rect 100076 37924 100082 37936
rect 103486 37924 103514 38168
rect 156046 38156 156052 38168
rect 156104 38156 156110 38208
rect 160738 38156 160744 38208
rect 160796 38196 160802 38208
rect 165982 38196 165988 38208
rect 160796 38168 165988 38196
rect 160796 38156 160802 38168
rect 165982 38156 165988 38168
rect 166040 38156 166046 38208
rect 201586 38156 201592 38208
rect 201644 38196 201650 38208
rect 247678 38196 247684 38208
rect 201644 38168 247684 38196
rect 201644 38156 201650 38168
rect 247678 38156 247684 38168
rect 247736 38156 247742 38208
rect 108298 38088 108304 38140
rect 108356 38128 108362 38140
rect 168834 38128 168840 38140
rect 108356 38100 168840 38128
rect 108356 38088 108362 38100
rect 168834 38088 168840 38100
rect 168892 38088 168898 38140
rect 169018 38088 169024 38140
rect 169076 38128 169082 38140
rect 178862 38128 178868 38140
rect 169076 38100 178868 38128
rect 169076 38088 169082 38100
rect 178862 38088 178868 38100
rect 178920 38088 178926 38140
rect 208762 38088 208768 38140
rect 208820 38128 208826 38140
rect 251818 38128 251824 38140
rect 208820 38100 251824 38128
rect 208820 38088 208826 38100
rect 251818 38088 251824 38100
rect 251876 38088 251882 38140
rect 104158 38020 104164 38072
rect 104216 38060 104222 38072
rect 164602 38060 164608 38072
rect 104216 38032 164608 38060
rect 104216 38020 104222 38032
rect 164602 38020 164608 38032
rect 164660 38020 164666 38072
rect 164878 38020 164884 38072
rect 164936 38060 164942 38072
rect 170306 38060 170312 38072
rect 164936 38032 170312 38060
rect 164936 38020 164942 38032
rect 170306 38020 170312 38032
rect 170364 38020 170370 38072
rect 175918 38020 175924 38072
rect 175976 38060 175982 38072
rect 188798 38060 188804 38072
rect 175976 38032 188804 38060
rect 175976 38020 175982 38032
rect 188798 38020 188804 38032
rect 188856 38020 188862 38072
rect 221550 38020 221556 38072
rect 221608 38060 221614 38072
rect 239490 38060 239496 38072
rect 221608 38032 239496 38060
rect 221608 38020 221614 38032
rect 239490 38020 239496 38032
rect 239548 38020 239554 38072
rect 104894 37952 104900 38004
rect 104952 37992 104958 38004
rect 106182 37992 106188 38004
rect 104952 37964 106188 37992
rect 104952 37952 104958 37964
rect 106182 37952 106188 37964
rect 106240 37952 106246 38004
rect 106274 37952 106280 38004
rect 106332 37992 106338 38004
rect 107562 37992 107568 38004
rect 106332 37964 107568 37992
rect 106332 37952 106338 37964
rect 107562 37952 107568 37964
rect 107620 37952 107626 38004
rect 115198 37952 115204 38004
rect 115256 37992 115262 38004
rect 177390 37992 177396 38004
rect 115256 37964 177396 37992
rect 115256 37952 115262 37964
rect 177390 37952 177396 37964
rect 177448 37952 177454 38004
rect 178678 37952 178684 38004
rect 178736 37992 178742 38004
rect 190270 37992 190276 38004
rect 178736 37964 190276 37992
rect 178736 37952 178742 37964
rect 190270 37952 190276 37964
rect 190328 37952 190334 38004
rect 205910 37952 205916 38004
rect 205968 37992 205974 38004
rect 375466 37992 375472 38004
rect 205968 37964 375472 37992
rect 205968 37952 205974 37964
rect 375466 37952 375472 37964
rect 375524 37952 375530 38004
rect 100076 37896 103514 37924
rect 100076 37884 100082 37896
rect 122098 37884 122104 37936
rect 122156 37924 122162 37936
rect 185946 37924 185952 37936
rect 122156 37896 185952 37924
rect 122156 37884 122162 37896
rect 185946 37884 185952 37896
rect 186004 37884 186010 37936
rect 217318 37884 217324 37936
rect 217376 37924 217382 37936
rect 382918 37924 382924 37936
rect 217376 37896 382924 37924
rect 217376 37884 217382 37896
rect 382918 37884 382924 37896
rect 382976 37884 382982 37936
rect 51718 37816 51724 37868
rect 51776 37856 51782 37868
rect 53466 37856 53472 37868
rect 51776 37828 53472 37856
rect 51776 37816 51782 37828
rect 53466 37816 53472 37828
rect 53524 37816 53530 37868
rect 57974 37816 57980 37868
rect 58032 37856 58038 37868
rect 59170 37856 59176 37868
rect 58032 37828 59176 37856
rect 58032 37816 58038 37828
rect 59170 37816 59176 37828
rect 59228 37816 59234 37868
rect 60734 37816 60740 37868
rect 60792 37856 60798 37868
rect 62022 37856 62028 37868
rect 60792 37828 62028 37856
rect 60792 37816 60798 37828
rect 62022 37816 62028 37828
rect 62080 37816 62086 37868
rect 149054 37816 149060 37868
rect 149112 37856 149118 37868
rect 150342 37856 150348 37868
rect 149112 37828 150348 37856
rect 149112 37816 149118 37828
rect 150342 37816 150348 37828
rect 150400 37816 150406 37868
rect 172606 37816 172612 37868
rect 172664 37856 172670 37868
rect 174538 37856 174544 37868
rect 172664 37828 174544 37856
rect 172664 37816 172670 37828
rect 174538 37816 174544 37828
rect 174596 37816 174602 37868
rect 203058 37816 203064 37868
rect 203116 37856 203122 37868
rect 371878 37856 371884 37868
rect 203116 37828 371884 37856
rect 203116 37816 203122 37828
rect 371878 37816 371884 37828
rect 371936 37816 371942 37868
rect 211614 37748 211620 37800
rect 211672 37788 211678 37800
rect 371326 37788 371332 37800
rect 211672 37760 371332 37788
rect 211672 37748 211678 37760
rect 371326 37748 371332 37760
rect 371384 37748 371390 37800
rect 55858 37680 55864 37732
rect 55916 37720 55922 37732
rect 63402 37720 63408 37732
rect 55916 37692 63408 37720
rect 55916 37680 55922 37692
rect 63402 37680 63408 37692
rect 63460 37680 63466 37732
rect 69658 37680 69664 37732
rect 69716 37720 69722 37732
rect 70578 37720 70584 37732
rect 69716 37692 70584 37720
rect 69716 37680 69722 37692
rect 70578 37680 70584 37692
rect 70636 37680 70642 37732
rect 113818 37680 113824 37732
rect 113876 37720 113882 37732
rect 114738 37720 114744 37732
rect 113876 37692 114744 37720
rect 113876 37680 113882 37692
rect 114738 37680 114744 37692
rect 114796 37680 114802 37732
rect 147674 37680 147680 37732
rect 147732 37720 147738 37732
rect 148870 37720 148876 37732
rect 147732 37692 148876 37720
rect 147732 37680 147738 37692
rect 148870 37680 148876 37692
rect 148928 37680 148934 37732
rect 174538 37680 174544 37732
rect 174596 37720 174602 37732
rect 180242 37720 180248 37732
rect 174596 37692 180248 37720
rect 174596 37680 174602 37692
rect 180242 37680 180248 37692
rect 180300 37680 180306 37732
rect 214466 37680 214472 37732
rect 214524 37720 214530 37732
rect 239674 37720 239680 37732
rect 214524 37692 239680 37720
rect 214524 37680 214530 37692
rect 239674 37680 239680 37692
rect 239732 37680 239738 37732
rect 218698 37612 218704 37664
rect 218756 37652 218762 37664
rect 239398 37652 239404 37664
rect 218756 37624 239404 37652
rect 218756 37612 218762 37624
rect 239398 37612 239404 37624
rect 239456 37612 239462 37664
rect 238662 37544 238668 37596
rect 238720 37584 238726 37596
rect 242986 37584 242992 37596
rect 238720 37556 242992 37584
rect 238720 37544 238726 37556
rect 242986 37544 242992 37556
rect 243044 37544 243050 37596
rect 48958 37476 48964 37528
rect 49016 37516 49022 37528
rect 51994 37516 52000 37528
rect 49016 37488 52000 37516
rect 49016 37476 49022 37488
rect 51994 37476 52000 37488
rect 52052 37476 52058 37528
rect 146938 37408 146944 37460
rect 146996 37448 147002 37460
rect 151722 37448 151728 37460
rect 146996 37420 151728 37448
rect 146996 37408 147002 37420
rect 151722 37408 151728 37420
rect 151780 37408 151786 37460
rect 54478 37272 54484 37324
rect 54536 37312 54542 37324
rect 57698 37312 57704 37324
rect 54536 37284 57704 37312
rect 54536 37272 54542 37284
rect 57698 37272 57704 37284
rect 57756 37272 57762 37324
rect 177298 37272 177304 37324
rect 177356 37312 177362 37324
rect 181714 37312 181720 37324
rect 177356 37284 181720 37312
rect 177356 37272 177362 37284
rect 181714 37272 181720 37284
rect 181772 37272 181778 37324
rect 19978 37136 19984 37188
rect 20036 37176 20042 37188
rect 54846 37176 54852 37188
rect 20036 37148 54852 37176
rect 20036 37136 20042 37148
rect 54846 37136 54852 37148
rect 54904 37136 54910 37188
rect 75178 37136 75184 37188
rect 75236 37176 75242 37188
rect 99006 37176 99012 37188
rect 75236 37148 99012 37176
rect 75236 37136 75242 37148
rect 99006 37136 99012 37148
rect 99064 37136 99070 37188
rect 8202 37068 8208 37120
rect 8260 37108 8266 37120
rect 49142 37108 49148 37120
rect 8260 37080 49148 37108
rect 8260 37068 8266 37080
rect 49142 37068 49148 37080
rect 49200 37068 49206 37120
rect 73798 37068 73804 37120
rect 73856 37108 73862 37120
rect 103330 37108 103336 37120
rect 73856 37080 103336 37108
rect 73856 37068 73862 37080
rect 103330 37068 103336 37080
rect 103388 37068 103394 37120
rect 32398 37000 32404 37052
rect 32456 37040 32462 37052
rect 76282 37040 76288 37052
rect 32456 37012 76288 37040
rect 32456 37000 32462 37012
rect 76282 37000 76288 37012
rect 76340 37000 76346 37052
rect 82078 37000 82084 37052
rect 82136 37040 82142 37052
rect 111886 37040 111892 37052
rect 82136 37012 111892 37040
rect 82136 37000 82142 37012
rect 111886 37000 111892 37012
rect 111944 37000 111950 37052
rect 34422 36932 34428 36984
rect 34480 36972 34486 36984
rect 80514 36972 80520 36984
rect 34480 36944 80520 36972
rect 34480 36932 34486 36944
rect 80514 36932 80520 36944
rect 80572 36932 80578 36984
rect 83458 36932 83464 36984
rect 83516 36972 83522 36984
rect 130378 36972 130384 36984
rect 83516 36944 130384 36972
rect 83516 36932 83522 36944
rect 130378 36932 130384 36944
rect 130436 36932 130442 36984
rect 15838 36864 15844 36916
rect 15896 36904 15902 36916
rect 43346 36904 43352 36916
rect 15896 36876 43352 36904
rect 15896 36864 15902 36876
rect 43346 36864 43352 36876
rect 43404 36864 43410 36916
rect 43438 36864 43444 36916
rect 43496 36904 43502 36916
rect 90542 36904 90548 36916
rect 43496 36876 90548 36904
rect 43496 36864 43502 36876
rect 90542 36864 90548 36876
rect 90600 36864 90606 36916
rect 95878 36864 95884 36916
rect 95936 36904 95942 36916
rect 113266 36904 113272 36916
rect 95936 36876 113272 36904
rect 95936 36864 95942 36876
rect 113266 36864 113272 36876
rect 113324 36864 113330 36916
rect 38562 36796 38568 36848
rect 38620 36836 38626 36848
rect 86218 36836 86224 36848
rect 38620 36808 86224 36836
rect 38620 36796 38626 36808
rect 86218 36796 86224 36808
rect 86276 36796 86282 36848
rect 91738 36796 91744 36848
rect 91796 36836 91802 36848
rect 116118 36836 116124 36848
rect 91796 36808 116124 36836
rect 91796 36796 91802 36808
rect 116118 36796 116124 36808
rect 116176 36796 116182 36848
rect 4062 36728 4068 36780
rect 4120 36768 4126 36780
rect 44910 36768 44916 36780
rect 4120 36740 44916 36768
rect 4120 36728 4126 36740
rect 44910 36728 44916 36740
rect 44968 36728 44974 36780
rect 53742 36728 53748 36780
rect 53800 36768 53806 36780
rect 104710 36768 104716 36780
rect 53800 36740 104716 36768
rect 53800 36728 53806 36740
rect 104710 36728 104716 36740
rect 104768 36728 104774 36780
rect 17862 36660 17868 36712
rect 17920 36700 17926 36712
rect 60550 36700 60556 36712
rect 17920 36672 60556 36700
rect 17920 36660 17926 36672
rect 60550 36660 60556 36672
rect 60608 36660 60614 36712
rect 68278 36660 68284 36712
rect 68336 36700 68342 36712
rect 118970 36700 118976 36712
rect 68336 36672 118976 36700
rect 68336 36660 68342 36672
rect 118970 36660 118976 36672
rect 119028 36660 119034 36712
rect 22002 36592 22008 36644
rect 22060 36632 22066 36644
rect 66254 36632 66260 36644
rect 22060 36604 66260 36632
rect 22060 36592 22066 36604
rect 66254 36592 66260 36604
rect 66312 36592 66318 36644
rect 71038 36592 71044 36644
rect 71096 36632 71102 36644
rect 123294 36632 123300 36644
rect 71096 36604 123300 36632
rect 71096 36592 71102 36604
rect 123294 36592 123300 36604
rect 123352 36592 123358 36644
rect 123478 36592 123484 36644
rect 123536 36632 123542 36644
rect 176010 36632 176016 36644
rect 123536 36604 176016 36632
rect 123536 36592 123542 36604
rect 176010 36592 176016 36604
rect 176068 36592 176074 36644
rect 2038 36524 2044 36576
rect 2096 36564 2102 36576
rect 40678 36564 40684 36576
rect 2096 36536 40684 36564
rect 2096 36524 2102 36536
rect 40678 36524 40684 36536
rect 40736 36524 40742 36576
rect 57882 36524 57888 36576
rect 57940 36564 57946 36576
rect 109034 36564 109040 36576
rect 57940 36536 109040 36564
rect 57940 36524 57946 36536
rect 109034 36524 109040 36536
rect 109092 36524 109098 36576
rect 119982 36524 119988 36576
rect 120040 36564 120046 36576
rect 184566 36564 184572 36576
rect 120040 36536 184572 36564
rect 120040 36524 120046 36536
rect 184566 36524 184572 36536
rect 184624 36524 184630 36576
rect 87598 35912 87604 35964
rect 87656 35952 87662 35964
rect 94774 35952 94780 35964
rect 87656 35924 94780 35952
rect 87656 35912 87662 35924
rect 94774 35912 94780 35924
rect 94832 35912 94838 35964
rect 126238 35912 126244 35964
rect 126296 35952 126302 35964
rect 134702 35952 134708 35964
rect 126296 35924 134708 35952
rect 126296 35912 126302 35924
rect 134702 35912 134708 35924
rect 134760 35912 134766 35964
rect 25498 35504 25504 35556
rect 25556 35544 25562 35556
rect 60734 35544 60740 35556
rect 25556 35516 60740 35544
rect 25556 35504 25562 35516
rect 60734 35504 60740 35516
rect 60792 35504 60798 35556
rect 35802 35436 35808 35488
rect 35860 35476 35866 35488
rect 81986 35476 81992 35488
rect 35860 35448 81992 35476
rect 35860 35436 35866 35448
rect 81986 35436 81992 35448
rect 82044 35436 82050 35488
rect 28902 35368 28908 35420
rect 28960 35408 28966 35420
rect 73430 35408 73436 35420
rect 28960 35380 73436 35408
rect 28960 35368 28966 35380
rect 73430 35368 73436 35380
rect 73488 35368 73494 35420
rect 77938 35368 77944 35420
rect 77996 35408 78002 35420
rect 126146 35408 126152 35420
rect 77996 35380 126152 35408
rect 77996 35368 78002 35380
rect 126146 35368 126152 35380
rect 126204 35368 126210 35420
rect 24118 35300 24124 35352
rect 24176 35340 24182 35352
rect 50614 35340 50620 35352
rect 24176 35312 50620 35340
rect 24176 35300 24182 35312
rect 50614 35300 50620 35312
rect 50672 35300 50678 35352
rect 50982 35300 50988 35352
rect 51040 35340 51046 35352
rect 99374 35340 99380 35352
rect 51040 35312 99380 35340
rect 51040 35300 51046 35312
rect 99374 35300 99380 35312
rect 99432 35300 99438 35352
rect 31662 35232 31668 35284
rect 31720 35272 31726 35284
rect 77662 35272 77668 35284
rect 31720 35244 77668 35272
rect 31720 35232 31726 35244
rect 77662 35232 77668 35244
rect 77720 35232 77726 35284
rect 86218 35232 86224 35284
rect 86276 35272 86282 35284
rect 138934 35272 138940 35284
rect 86276 35244 138940 35272
rect 86276 35232 86282 35244
rect 138934 35232 138940 35244
rect 138992 35232 138998 35284
rect 13722 35164 13728 35216
rect 13780 35204 13786 35216
rect 55214 35204 55220 35216
rect 13780 35176 55220 35204
rect 13780 35164 13786 35176
rect 55214 35164 55220 35176
rect 55272 35164 55278 35216
rect 64782 35164 64788 35216
rect 64840 35204 64846 35216
rect 117590 35204 117596 35216
rect 64840 35176 117596 35204
rect 64840 35164 64846 35176
rect 117590 35164 117596 35176
rect 117648 35164 117654 35216
rect 117958 34484 117964 34536
rect 118016 34524 118022 34536
rect 121822 34524 121828 34536
rect 118016 34496 121828 34524
rect 118016 34484 118022 34496
rect 121822 34484 121828 34496
rect 121880 34484 121886 34536
rect 266998 33056 267004 33108
rect 267056 33096 267062 33108
rect 580166 33096 580172 33108
rect 267056 33068 580172 33096
rect 267056 33056 267062 33068
rect 580166 33056 580172 33068
rect 580224 33056 580230 33108
rect 2774 32784 2780 32836
rect 2832 32824 2838 32836
rect 6178 32824 6184 32836
rect 2832 32796 6184 32824
rect 2832 32784 2838 32796
rect 6178 32784 6184 32796
rect 6236 32784 6242 32836
rect 6270 32376 6276 32428
rect 6328 32416 6334 32428
rect 46290 32416 46296 32428
rect 6328 32388 46296 32416
rect 6328 32376 6334 32388
rect 46290 32376 46296 32388
rect 46348 32376 46354 32428
rect 111702 29588 111708 29640
rect 111760 29628 111766 29640
rect 172606 29628 172612 29640
rect 111760 29600 172612 29628
rect 111760 29588 111766 29600
rect 172606 29588 172612 29600
rect 172664 29588 172670 29640
rect 3418 20612 3424 20664
rect 3476 20652 3482 20664
rect 14458 20652 14464 20664
rect 3476 20624 14464 20652
rect 3476 20612 3482 20624
rect 14458 20612 14464 20624
rect 14516 20612 14522 20664
rect 276658 20612 276664 20664
rect 276716 20652 276722 20664
rect 580166 20652 580172 20664
rect 276716 20624 580172 20652
rect 276716 20612 276722 20624
rect 580166 20612 580172 20624
rect 580224 20612 580230 20664
rect 88242 8916 88248 8968
rect 88300 8956 88306 8968
rect 132494 8956 132500 8968
rect 88300 8928 132500 8956
rect 88300 8916 88306 8928
rect 132494 8916 132500 8928
rect 132552 8916 132558 8968
rect 24762 7556 24768 7608
rect 24820 7596 24826 7608
rect 67634 7596 67640 7608
rect 24820 7568 67640 7596
rect 24820 7556 24826 7568
rect 67634 7556 67640 7568
rect 67692 7556 67698 7608
rect 95326 7556 95332 7608
rect 95384 7596 95390 7608
rect 153194 7596 153200 7608
rect 95384 7568 153200 7596
rect 95384 7556 95390 7568
rect 153194 7556 153200 7568
rect 153252 7556 153258 7608
rect 3418 6808 3424 6860
rect 3476 6848 3482 6860
rect 10318 6848 10324 6860
rect 3476 6820 10324 6848
rect 3476 6808 3482 6820
rect 10318 6808 10324 6820
rect 10376 6808 10382 6860
rect 85206 6604 85212 6656
rect 85264 6644 85270 6656
rect 136634 6644 136640 6656
rect 85264 6616 136640 6644
rect 85264 6604 85270 6616
rect 136634 6604 136640 6616
rect 136692 6604 136698 6656
rect 61654 6536 61660 6588
rect 61712 6576 61718 6588
rect 110414 6576 110420 6588
rect 61712 6548 110420 6576
rect 61712 6536 61718 6548
rect 110414 6536 110420 6548
rect 110472 6536 110478 6588
rect 115290 6536 115296 6588
rect 115348 6576 115354 6588
rect 169018 6576 169024 6588
rect 115348 6548 169024 6576
rect 115348 6536 115354 6548
rect 169018 6536 169024 6548
rect 169076 6536 169082 6588
rect 108114 6468 108120 6520
rect 108172 6508 108178 6520
rect 164878 6508 164884 6520
rect 108172 6480 164884 6508
rect 108172 6468 108178 6480
rect 164878 6468 164884 6480
rect 164936 6468 164942 6520
rect 104526 6400 104532 6452
rect 104584 6440 104590 6452
rect 160738 6440 160744 6452
rect 104584 6412 160744 6440
rect 104584 6400 104590 6412
rect 160738 6400 160744 6412
rect 160796 6400 160802 6452
rect 51350 6332 51356 6384
rect 51408 6372 51414 6384
rect 100754 6372 100760 6384
rect 51408 6344 100760 6372
rect 51408 6332 51414 6344
rect 100754 6332 100760 6344
rect 100812 6332 100818 6384
rect 101030 6332 101036 6384
rect 101088 6372 101094 6384
rect 161474 6372 161480 6384
rect 101088 6344 161480 6372
rect 101088 6332 101094 6344
rect 161474 6332 161480 6344
rect 161532 6332 161538 6384
rect 47854 6264 47860 6316
rect 47912 6304 47918 6316
rect 96614 6304 96620 6316
rect 47912 6276 96620 6304
rect 47912 6264 47918 6276
rect 96614 6264 96620 6276
rect 96672 6264 96678 6316
rect 97442 6264 97448 6316
rect 97500 6304 97506 6316
rect 157334 6304 157340 6316
rect 97500 6276 157340 6304
rect 97500 6264 97506 6276
rect 157334 6264 157340 6276
rect 157392 6264 157398 6316
rect 54938 6196 54944 6248
rect 54996 6236 55002 6248
rect 104894 6236 104900 6248
rect 54996 6208 104900 6236
rect 54996 6196 55002 6208
rect 104894 6196 104900 6208
rect 104952 6196 104958 6248
rect 118786 6196 118792 6248
rect 118844 6236 118850 6248
rect 182174 6236 182180 6248
rect 118844 6208 182180 6236
rect 118844 6196 118850 6208
rect 182174 6196 182180 6208
rect 182232 6196 182238 6248
rect 62022 6128 62028 6180
rect 62080 6168 62086 6180
rect 113818 6168 113824 6180
rect 62080 6140 113824 6168
rect 62080 6128 62086 6140
rect 113818 6128 113824 6140
rect 113876 6128 113882 6180
rect 122282 6128 122288 6180
rect 122340 6168 122346 6180
rect 186314 6168 186320 6180
rect 122340 6140 186320 6168
rect 122340 6128 122346 6140
rect 186314 6128 186320 6140
rect 186372 6128 186378 6180
rect 76190 5448 76196 5500
rect 76248 5488 76254 5500
rect 131114 5488 131120 5500
rect 76248 5460 131120 5488
rect 76248 5448 76254 5460
rect 131114 5448 131120 5460
rect 131172 5448 131178 5500
rect 72602 5380 72608 5432
rect 72660 5420 72666 5432
rect 126974 5420 126980 5432
rect 72660 5392 126980 5420
rect 72660 5380 72666 5392
rect 126974 5380 126980 5392
rect 127032 5380 127038 5432
rect 70302 5312 70308 5364
rect 70360 5352 70366 5364
rect 124214 5352 124220 5364
rect 70360 5324 124220 5352
rect 70360 5312 70366 5324
rect 124214 5312 124220 5324
rect 124272 5312 124278 5364
rect 79686 5244 79692 5296
rect 79744 5284 79750 5296
rect 135254 5284 135260 5296
rect 79744 5256 135260 5284
rect 79744 5244 79750 5256
rect 135254 5244 135260 5256
rect 135312 5244 135318 5296
rect 83274 5176 83280 5228
rect 83332 5216 83338 5228
rect 139394 5216 139400 5228
rect 83332 5188 139400 5216
rect 83332 5176 83338 5188
rect 139394 5176 139400 5188
rect 139452 5176 139458 5228
rect 86862 5108 86868 5160
rect 86920 5148 86926 5160
rect 143534 5148 143540 5160
rect 86920 5120 143540 5148
rect 86920 5108 86926 5120
rect 143534 5108 143540 5120
rect 143592 5108 143598 5160
rect 90450 5040 90456 5092
rect 90508 5080 90514 5092
rect 147674 5080 147680 5092
rect 90508 5052 147680 5080
rect 90508 5040 90514 5052
rect 147674 5040 147680 5052
rect 147732 5040 147738 5092
rect 28994 4972 29000 5024
rect 29052 5012 29058 5024
rect 71774 5012 71780 5024
rect 29052 4984 71780 5012
rect 29052 4972 29058 4984
rect 71774 4972 71780 4984
rect 71832 4972 71838 5024
rect 87966 4972 87972 5024
rect 88024 5012 88030 5024
rect 144914 5012 144920 5024
rect 88024 4984 144920 5012
rect 88024 4972 88030 4984
rect 144914 4972 144920 4984
rect 144972 4972 144978 5024
rect 40678 4904 40684 4956
rect 40736 4944 40742 4956
rect 88334 4944 88340 4956
rect 40736 4916 88340 4944
rect 40736 4904 40742 4916
rect 88334 4904 88340 4916
rect 88392 4904 88398 4956
rect 102226 4904 102232 4956
rect 102284 4944 102290 4956
rect 162854 4944 162860 4956
rect 102284 4916 162860 4944
rect 102284 4904 102290 4916
rect 162854 4904 162860 4916
rect 162912 4904 162918 4956
rect 37182 4836 37188 4888
rect 37240 4876 37246 4888
rect 84194 4876 84200 4888
rect 37240 4848 84200 4876
rect 37240 4836 37246 4848
rect 84194 4836 84200 4848
rect 84252 4836 84258 4888
rect 95142 4836 95148 4888
rect 95200 4876 95206 4888
rect 154574 4876 154580 4888
rect 95200 4848 154580 4876
rect 95200 4836 95206 4848
rect 154574 4836 154580 4848
rect 154632 4836 154638 4888
rect 9950 4768 9956 4820
rect 10008 4808 10014 4820
rect 48958 4808 48964 4820
rect 10008 4780 48964 4808
rect 10008 4768 10014 4780
rect 48958 4768 48964 4780
rect 49016 4768 49022 4820
rect 56042 4768 56048 4820
rect 56100 4808 56106 4820
rect 106274 4808 106280 4820
rect 56100 4780 106280 4808
rect 56100 4768 56106 4780
rect 106274 4768 106280 4780
rect 106332 4768 106338 4820
rect 109310 4768 109316 4820
rect 109368 4808 109374 4820
rect 171134 4808 171140 4820
rect 109368 4780 171140 4808
rect 109368 4768 109374 4780
rect 171134 4768 171140 4780
rect 171192 4768 171198 4820
rect 73798 4700 73804 4752
rect 73856 4740 73862 4752
rect 128354 4740 128360 4752
rect 73856 4712 128360 4740
rect 73856 4700 73862 4712
rect 128354 4700 128360 4712
rect 128412 4700 128418 4752
rect 66714 4632 66720 4684
rect 66772 4672 66778 4684
rect 120074 4672 120080 4684
rect 66772 4644 120080 4672
rect 66772 4632 66778 4644
rect 120074 4632 120080 4644
rect 120132 4632 120138 4684
rect 43070 4088 43076 4140
rect 43128 4128 43134 4140
rect 79318 4128 79324 4140
rect 43128 4100 79324 4128
rect 43128 4088 43134 4100
rect 79318 4088 79324 4100
rect 79376 4088 79382 4140
rect 103330 4088 103336 4140
rect 103388 4128 103394 4140
rect 104158 4128 104164 4140
rect 103388 4100 104164 4128
rect 103388 4088 103394 4100
rect 104158 4088 104164 4100
rect 104216 4088 104222 4140
rect 123478 4088 123484 4140
rect 123536 4128 123542 4140
rect 175918 4128 175924 4140
rect 123536 4100 175924 4128
rect 123536 4088 123542 4100
rect 175918 4088 175924 4100
rect 175976 4088 175982 4140
rect 19426 4020 19432 4072
rect 19484 4060 19490 4072
rect 50341 4063 50399 4069
rect 50341 4060 50353 4063
rect 19484 4032 50353 4060
rect 19484 4020 19490 4032
rect 50341 4029 50353 4032
rect 50387 4029 50399 4063
rect 50341 4023 50399 4029
rect 50433 4063 50491 4069
rect 50433 4029 50445 4063
rect 50479 4060 50491 4063
rect 54478 4060 54484 4072
rect 50479 4032 54484 4060
rect 50479 4029 50491 4032
rect 50433 4023 50491 4029
rect 54478 4020 54484 4032
rect 54536 4020 54542 4072
rect 91738 4060 91744 4072
rect 64846 4032 91744 4060
rect 24210 3952 24216 4004
rect 24268 3992 24274 4004
rect 59998 3992 60004 4004
rect 24268 3964 60004 3992
rect 24268 3952 24274 3964
rect 59998 3952 60004 3964
rect 60056 3952 60062 4004
rect 63218 3952 63224 4004
rect 63276 3992 63282 4004
rect 64846 3992 64874 4032
rect 91738 4020 91744 4032
rect 91796 4020 91802 4072
rect 92750 4020 92756 4072
rect 92808 4060 92814 4072
rect 146938 4060 146944 4072
rect 92808 4032 146944 4060
rect 92808 4020 92814 4032
rect 146938 4020 146944 4032
rect 146996 4020 147002 4072
rect 63276 3964 64874 3992
rect 63276 3952 63282 3964
rect 67910 3952 67916 4004
rect 67968 3992 67974 4004
rect 117958 3992 117964 4004
rect 67968 3964 117964 3992
rect 67968 3952 67974 3964
rect 117958 3952 117964 3964
rect 118016 3952 118022 4004
rect 124674 3952 124680 4004
rect 124732 3992 124738 4004
rect 178678 3992 178684 4004
rect 124732 3964 178684 3992
rect 124732 3952 124738 3964
rect 178678 3952 178684 3964
rect 178736 3952 178742 4004
rect 11146 3884 11152 3936
rect 11204 3924 11210 3936
rect 51718 3924 51724 3936
rect 11204 3896 51724 3924
rect 11204 3884 11210 3896
rect 51718 3884 51724 3896
rect 51776 3884 51782 3936
rect 52546 3884 52552 3936
rect 52604 3924 52610 3936
rect 73706 3924 73712 3936
rect 52604 3896 73712 3924
rect 52604 3884 52610 3896
rect 73706 3884 73712 3896
rect 73764 3884 73770 3936
rect 85666 3884 85672 3936
rect 85724 3924 85730 3936
rect 142154 3924 142160 3936
rect 85724 3896 142160 3924
rect 85724 3884 85730 3896
rect 142154 3884 142160 3896
rect 142212 3884 142218 3936
rect 14734 3816 14740 3868
rect 14792 3856 14798 3868
rect 50249 3859 50307 3865
rect 50249 3856 50261 3859
rect 14792 3828 50261 3856
rect 14792 3816 14798 3828
rect 50249 3825 50261 3828
rect 50295 3825 50307 3859
rect 50249 3819 50307 3825
rect 50341 3859 50399 3865
rect 50341 3825 50353 3859
rect 50387 3856 50399 3859
rect 55858 3856 55864 3868
rect 50387 3828 55864 3856
rect 50387 3825 50399 3828
rect 50341 3819 50399 3825
rect 55858 3816 55864 3828
rect 55916 3816 55922 3868
rect 59630 3816 59636 3868
rect 59688 3856 59694 3868
rect 81986 3856 81992 3868
rect 59688 3828 81992 3856
rect 59688 3816 59694 3828
rect 81986 3816 81992 3828
rect 82044 3816 82050 3868
rect 82078 3816 82084 3868
rect 82136 3856 82142 3868
rect 82136 3828 84194 3856
rect 82136 3816 82142 3828
rect 6454 3748 6460 3800
rect 6512 3788 6518 3800
rect 46934 3788 46940 3800
rect 6512 3760 46940 3788
rect 6512 3748 6518 3760
rect 46934 3748 46940 3760
rect 46992 3748 46998 3800
rect 48958 3748 48964 3800
rect 49016 3788 49022 3800
rect 69661 3791 69719 3797
rect 69661 3788 69673 3791
rect 49016 3760 69673 3788
rect 49016 3748 49022 3760
rect 69661 3757 69673 3760
rect 69707 3757 69719 3791
rect 84166 3788 84194 3828
rect 84470 3816 84476 3868
rect 84528 3856 84534 3868
rect 140774 3856 140780 3868
rect 84528 3828 140780 3856
rect 84528 3816 84534 3828
rect 140774 3816 140780 3828
rect 140832 3816 140838 3868
rect 86218 3788 86224 3800
rect 84166 3760 86224 3788
rect 69661 3751 69719 3757
rect 86218 3748 86224 3760
rect 86276 3748 86282 3800
rect 91554 3748 91560 3800
rect 91612 3788 91618 3800
rect 149054 3788 149060 3800
rect 91612 3760 149060 3788
rect 91612 3748 91618 3760
rect 149054 3748 149060 3760
rect 149112 3748 149118 3800
rect 15930 3680 15936 3732
rect 15988 3720 15994 3732
rect 57974 3720 57980 3732
rect 15988 3692 57980 3720
rect 15988 3680 15994 3692
rect 57974 3680 57980 3692
rect 58032 3680 58038 3732
rect 60826 3680 60832 3732
rect 60884 3720 60890 3732
rect 95878 3720 95884 3732
rect 60884 3692 95884 3720
rect 60884 3680 60890 3692
rect 95878 3680 95884 3692
rect 95936 3680 95942 3732
rect 117590 3680 117596 3732
rect 117648 3720 117654 3732
rect 122285 3723 122343 3729
rect 117648 3692 122236 3720
rect 117648 3680 117654 3692
rect 30098 3612 30104 3664
rect 30156 3652 30162 3664
rect 32398 3652 32404 3664
rect 30156 3624 32404 3652
rect 30156 3612 30162 3624
rect 32398 3612 32404 3624
rect 32456 3612 32462 3664
rect 45462 3612 45468 3664
rect 45520 3652 45526 3664
rect 87598 3652 87604 3664
rect 45520 3624 87604 3652
rect 45520 3612 45526 3624
rect 87598 3612 87604 3624
rect 87656 3612 87662 3664
rect 114002 3612 114008 3664
rect 114060 3652 114066 3664
rect 115198 3652 115204 3664
rect 114060 3624 115204 3652
rect 114060 3612 114066 3624
rect 115198 3612 115204 3624
rect 115256 3612 115262 3664
rect 121086 3612 121092 3664
rect 121144 3652 121150 3664
rect 122098 3652 122104 3664
rect 121144 3624 122104 3652
rect 121144 3612 121150 3624
rect 122098 3612 122104 3624
rect 122156 3612 122162 3664
rect 122208 3652 122236 3692
rect 122285 3689 122297 3723
rect 122331 3720 122343 3723
rect 174538 3720 174544 3732
rect 122331 3692 174544 3720
rect 122331 3689 122343 3692
rect 122285 3683 122343 3689
rect 174538 3680 174544 3692
rect 174596 3680 174602 3732
rect 177298 3652 177304 3664
rect 122208 3624 177304 3652
rect 177298 3612 177304 3624
rect 177356 3612 177362 3664
rect 1670 3544 1676 3596
rect 1728 3584 1734 3596
rect 10318 3584 10324 3596
rect 1728 3556 10324 3584
rect 1728 3544 1734 3556
rect 10318 3544 10324 3556
rect 10376 3544 10382 3596
rect 12342 3544 12348 3596
rect 12400 3584 12406 3596
rect 19978 3584 19984 3596
rect 12400 3556 19984 3584
rect 12400 3544 12406 3556
rect 19978 3544 19984 3556
rect 20036 3544 20042 3596
rect 25314 3544 25320 3596
rect 25372 3584 25378 3596
rect 69658 3584 69664 3596
rect 25372 3556 69664 3584
rect 25372 3544 25378 3556
rect 69658 3544 69664 3556
rect 69716 3544 69722 3596
rect 74994 3544 75000 3596
rect 75052 3584 75058 3596
rect 83458 3584 83464 3596
rect 75052 3556 83464 3584
rect 75052 3544 75058 3556
rect 83458 3544 83464 3556
rect 83516 3544 83522 3596
rect 98638 3544 98644 3596
rect 98696 3584 98702 3596
rect 158714 3584 158720 3596
rect 98696 3556 158720 3584
rect 98696 3544 98702 3556
rect 158714 3544 158720 3556
rect 158772 3544 158778 3596
rect 193122 3544 193128 3596
rect 193180 3584 193186 3596
rect 582190 3584 582196 3596
rect 193180 3556 582196 3584
rect 193180 3544 193186 3556
rect 582190 3544 582196 3556
rect 582248 3544 582254 3596
rect 5258 3476 5264 3528
rect 5316 3516 5322 3528
rect 6270 3516 6276 3528
rect 5316 3488 6276 3516
rect 5316 3476 5322 3488
rect 6270 3476 6276 3488
rect 6328 3476 6334 3528
rect 7650 3476 7656 3528
rect 7708 3516 7714 3528
rect 8202 3516 8208 3528
rect 7708 3488 8208 3516
rect 7708 3476 7714 3488
rect 8202 3476 8208 3488
rect 8260 3476 8266 3528
rect 17034 3476 17040 3528
rect 17092 3516 17098 3528
rect 17862 3516 17868 3528
rect 17092 3488 17868 3516
rect 17092 3476 17098 3488
rect 17862 3476 17868 3488
rect 17920 3476 17926 3528
rect 23014 3476 23020 3528
rect 23072 3516 23078 3528
rect 24762 3516 24768 3528
rect 23072 3488 24768 3516
rect 23072 3476 23078 3488
rect 24762 3476 24768 3488
rect 24820 3476 24826 3528
rect 64874 3516 64880 3528
rect 26206 3488 64880 3516
rect 2866 3408 2872 3460
rect 2924 3448 2930 3460
rect 15838 3448 15844 3460
rect 2924 3420 15844 3448
rect 2924 3408 2930 3420
rect 15838 3408 15844 3420
rect 15896 3408 15902 3460
rect 20622 3408 20628 3460
rect 20680 3448 20686 3460
rect 26206 3448 26234 3488
rect 64874 3476 64880 3488
rect 64932 3476 64938 3528
rect 65518 3476 65524 3528
rect 65576 3516 65582 3528
rect 68278 3516 68284 3528
rect 65576 3488 68284 3516
rect 65576 3476 65582 3488
rect 68278 3476 68284 3488
rect 68336 3476 68342 3528
rect 69106 3476 69112 3528
rect 69164 3516 69170 3528
rect 71038 3516 71044 3528
rect 69164 3488 71044 3516
rect 69164 3476 69170 3488
rect 71038 3476 71044 3488
rect 71096 3476 71102 3528
rect 77386 3476 77392 3528
rect 77444 3516 77450 3528
rect 88242 3516 88248 3528
rect 77444 3488 88248 3516
rect 77444 3476 77450 3488
rect 88242 3476 88248 3488
rect 88300 3476 88306 3528
rect 89162 3476 89168 3528
rect 89220 3516 89226 3528
rect 90358 3516 90364 3528
rect 89220 3488 90364 3516
rect 89220 3476 89226 3488
rect 90358 3476 90364 3488
rect 90416 3476 90422 3528
rect 93946 3476 93952 3528
rect 94004 3516 94010 3528
rect 95326 3516 95332 3528
rect 94004 3488 95332 3516
rect 94004 3476 94010 3488
rect 95326 3476 95332 3488
rect 95384 3476 95390 3528
rect 106918 3476 106924 3528
rect 106976 3516 106982 3528
rect 108298 3516 108304 3528
rect 106976 3488 108304 3516
rect 106976 3476 106982 3488
rect 108298 3476 108304 3488
rect 108356 3476 108362 3528
rect 110506 3476 110512 3528
rect 110564 3516 110570 3528
rect 172514 3516 172520 3528
rect 110564 3488 172520 3516
rect 110564 3476 110570 3488
rect 172514 3476 172520 3488
rect 172572 3476 172578 3528
rect 194502 3476 194508 3528
rect 194560 3516 194566 3528
rect 583386 3516 583392 3528
rect 194560 3488 583392 3516
rect 194560 3476 194566 3488
rect 583386 3476 583392 3488
rect 583444 3476 583450 3528
rect 20680 3420 26234 3448
rect 20680 3408 20686 3420
rect 27706 3408 27712 3460
rect 27764 3448 27770 3460
rect 28902 3448 28908 3460
rect 27764 3420 28908 3448
rect 27764 3408 27770 3420
rect 28902 3408 28908 3420
rect 28960 3408 28966 3460
rect 33594 3408 33600 3460
rect 33652 3448 33658 3460
rect 34422 3448 34428 3460
rect 33652 3420 34428 3448
rect 33652 3408 33658 3420
rect 34422 3408 34428 3420
rect 34480 3408 34486 3460
rect 34790 3408 34796 3460
rect 34848 3448 34854 3460
rect 35802 3448 35808 3460
rect 34848 3420 35808 3448
rect 34848 3408 34854 3420
rect 35802 3408 35808 3420
rect 35860 3408 35866 3460
rect 35986 3408 35992 3460
rect 36044 3448 36050 3460
rect 37090 3448 37096 3460
rect 36044 3420 37096 3448
rect 36044 3408 36050 3420
rect 37090 3408 37096 3420
rect 37148 3408 37154 3460
rect 41874 3408 41880 3460
rect 41932 3448 41938 3460
rect 43438 3448 43444 3460
rect 41932 3420 43444 3448
rect 41932 3408 41938 3420
rect 43438 3408 43444 3420
rect 43496 3408 43502 3460
rect 44266 3408 44272 3460
rect 44324 3448 44330 3460
rect 92474 3448 92480 3460
rect 44324 3420 92480 3448
rect 44324 3408 44330 3420
rect 92474 3408 92480 3420
rect 92532 3408 92538 3460
rect 105722 3408 105728 3460
rect 105780 3448 105786 3460
rect 166994 3448 167000 3460
rect 105780 3420 167000 3448
rect 105780 3408 105786 3420
rect 166994 3408 167000 3420
rect 167052 3408 167058 3460
rect 191742 3408 191748 3460
rect 191800 3448 191806 3460
rect 580994 3448 581000 3460
rect 191800 3420 581000 3448
rect 191800 3408 191806 3420
rect 580994 3408 581000 3420
rect 581052 3408 581058 3460
rect 566 3340 572 3392
rect 624 3380 630 3392
rect 2038 3380 2044 3392
rect 624 3352 2044 3380
rect 624 3340 630 3352
rect 2038 3340 2044 3352
rect 2096 3340 2102 3392
rect 8754 3340 8760 3392
rect 8812 3380 8818 3392
rect 24118 3380 24124 3392
rect 8812 3352 24124 3380
rect 8812 3340 8818 3352
rect 24118 3340 24124 3352
rect 24176 3340 24182 3392
rect 32398 3340 32404 3392
rect 32456 3380 32462 3392
rect 66898 3380 66904 3392
rect 32456 3352 66904 3380
rect 32456 3340 32462 3352
rect 66898 3340 66904 3352
rect 66956 3340 66962 3392
rect 71498 3340 71504 3392
rect 71556 3380 71562 3392
rect 77938 3380 77944 3392
rect 71556 3352 77944 3380
rect 71556 3340 71562 3352
rect 77938 3340 77944 3352
rect 77996 3340 78002 3392
rect 80882 3340 80888 3392
rect 80940 3380 80946 3392
rect 85206 3380 85212 3392
rect 80940 3352 85212 3380
rect 80940 3340 80946 3352
rect 85206 3340 85212 3352
rect 85264 3340 85270 3392
rect 99834 3340 99840 3392
rect 99892 3380 99898 3392
rect 151078 3380 151084 3392
rect 99892 3352 151084 3380
rect 99892 3340 99898 3352
rect 151078 3340 151084 3352
rect 151136 3340 151142 3392
rect 28902 3272 28908 3324
rect 28960 3312 28966 3324
rect 28960 3284 45554 3312
rect 28960 3272 28966 3284
rect 45526 3244 45554 3284
rect 50154 3272 50160 3324
rect 50212 3312 50218 3324
rect 50982 3312 50988 3324
rect 50212 3284 50988 3312
rect 50212 3272 50218 3284
rect 50982 3272 50988 3284
rect 51040 3272 51046 3324
rect 57238 3272 57244 3324
rect 57296 3312 57302 3324
rect 57882 3312 57888 3324
rect 57296 3284 57888 3312
rect 57296 3272 57302 3284
rect 57882 3272 57888 3284
rect 57940 3272 57946 3324
rect 58434 3272 58440 3324
rect 58492 3312 58498 3324
rect 61654 3312 61660 3324
rect 58492 3284 61660 3312
rect 58492 3272 58498 3284
rect 61654 3272 61660 3284
rect 61712 3272 61718 3324
rect 64322 3272 64328 3324
rect 64380 3312 64386 3324
rect 64782 3312 64788 3324
rect 64380 3284 64788 3312
rect 64380 3272 64386 3284
rect 64782 3272 64788 3284
rect 64840 3272 64846 3324
rect 69661 3315 69719 3321
rect 69661 3281 69673 3315
rect 69707 3312 69719 3315
rect 75178 3312 75184 3324
rect 69707 3284 75184 3312
rect 69707 3281 69719 3284
rect 69661 3275 69719 3281
rect 75178 3272 75184 3284
rect 75236 3272 75242 3324
rect 78582 3272 78588 3324
rect 78640 3312 78646 3324
rect 126238 3312 126244 3324
rect 78640 3284 126244 3312
rect 78640 3272 78646 3284
rect 126238 3272 126244 3284
rect 126296 3272 126302 3324
rect 61378 3244 61384 3256
rect 45526 3216 61384 3244
rect 61378 3204 61384 3216
rect 61436 3204 61442 3256
rect 112806 3204 112812 3256
rect 112864 3244 112870 3256
rect 123386 3244 123392 3256
rect 112864 3216 123392 3244
rect 112864 3204 112870 3216
rect 123386 3204 123392 3216
rect 123444 3204 123450 3256
rect 96246 3136 96252 3188
rect 96304 3176 96310 3188
rect 100018 3176 100024 3188
rect 96304 3148 100024 3176
rect 96304 3136 96310 3148
rect 100018 3136 100024 3148
rect 100076 3136 100082 3188
rect 116394 3136 116400 3188
rect 116452 3176 116458 3188
rect 122285 3179 122343 3185
rect 122285 3176 122297 3179
rect 116452 3148 122297 3176
rect 116452 3136 116458 3148
rect 122285 3145 122297 3148
rect 122331 3145 122343 3179
rect 122285 3139 122343 3145
rect 18230 2864 18236 2916
rect 18288 2904 18294 2916
rect 25498 2904 25504 2916
rect 18288 2876 25504 2904
rect 18288 2864 18294 2876
rect 25498 2864 25504 2876
rect 25556 2864 25562 2916
rect 26510 2796 26516 2848
rect 26568 2836 26574 2848
rect 28994 2836 29000 2848
rect 26568 2808 29000 2836
rect 26568 2796 26574 2808
rect 28994 2796 29000 2808
rect 29052 2796 29058 2848
<< via1 >>
rect 201500 702992 201552 703044
rect 202788 702992 202840 703044
rect 333244 700612 333296 700664
rect 364984 700612 365036 700664
rect 327724 700544 327776 700596
rect 429844 700544 429896 700596
rect 330484 700476 330536 700528
rect 462320 700476 462372 700528
rect 211804 700408 211856 700460
rect 348792 700408 348844 700460
rect 105452 700340 105504 700392
rect 106188 700340 106240 700392
rect 170312 700340 170364 700392
rect 178040 700340 178092 700392
rect 193864 700340 193916 700392
rect 332508 700340 332560 700392
rect 334624 700340 334676 700392
rect 397460 700340 397512 700392
rect 480904 700340 480956 700392
rect 494796 700340 494848 700392
rect 39856 700272 39908 700324
rect 89168 700272 89220 700324
rect 137836 700272 137888 700324
rect 176660 700272 176712 700324
rect 262864 700272 262916 700324
rect 413652 700272 413704 700324
rect 479524 700272 479576 700324
rect 559656 700272 559708 700324
rect 24308 699660 24360 699712
rect 24768 699660 24820 699712
rect 39764 699660 39816 699712
rect 40500 699660 40552 699712
rect 71780 699660 71832 699712
rect 72976 699660 73028 699712
rect 266360 697552 266412 697604
rect 267648 697552 267700 697604
rect 191104 696940 191156 696992
rect 580172 696940 580224 696992
rect 2780 683612 2832 683664
rect 6184 683612 6236 683664
rect 207664 683136 207716 683188
rect 580172 683136 580224 683188
rect 182824 670692 182876 670744
rect 580172 670692 580224 670744
rect 3516 656888 3568 656940
rect 15844 656888 15896 656940
rect 189724 643084 189776 643136
rect 580172 643084 580224 643136
rect 3516 632068 3568 632120
rect 35164 632068 35216 632120
rect 180064 616836 180116 616888
rect 580172 616836 580224 616888
rect 3332 605820 3384 605872
rect 17224 605820 17276 605872
rect 258724 590656 258776 590708
rect 580172 590656 580224 590708
rect 3332 579640 3384 579692
rect 31024 579640 31076 579692
rect 204904 576852 204956 576904
rect 580172 576852 580224 576904
rect 545764 563048 545816 563100
rect 580172 563048 580224 563100
rect 3332 553392 3384 553444
rect 28264 553392 28316 553444
rect 186964 536800 187016 536852
rect 579896 536800 579948 536852
rect 3332 527144 3384 527196
rect 10324 527144 10376 527196
rect 196624 524424 196676 524476
rect 580172 524424 580224 524476
rect 3332 514768 3384 514820
rect 32404 514768 32456 514820
rect 255964 510620 256016 510672
rect 580172 510620 580224 510672
rect 2872 500964 2924 501016
rect 33784 500964 33836 501016
rect 185584 484372 185636 484424
rect 580172 484372 580224 484424
rect 3332 474716 3384 474768
rect 13084 474716 13136 474768
rect 153200 473968 153252 474020
rect 176752 473968 176804 474020
rect 3332 462340 3384 462392
rect 21364 462340 21416 462392
rect 178684 456764 178736 456816
rect 580172 456764 580224 456816
rect 3332 448536 3384 448588
rect 19984 448536 20036 448588
rect 39672 425688 39724 425740
rect 71780 425688 71832 425740
rect 106188 425688 106240 425740
rect 176844 425688 176896 425740
rect 3148 422288 3200 422340
rect 25504 422288 25556 422340
rect 486424 418140 486476 418192
rect 580172 418140 580224 418192
rect 483664 404336 483716 404388
rect 580172 404336 580224 404388
rect 3332 397468 3384 397520
rect 21456 397468 21508 397520
rect 261484 376728 261536 376780
rect 337660 376728 337712 376780
rect 254584 375368 254636 375420
rect 337752 375368 337804 375420
rect 251824 372648 251876 372700
rect 337476 372648 337528 372700
rect 198648 372580 198700 372632
rect 337660 372580 337712 372632
rect 3332 371220 3384 371272
rect 14464 371220 14516 371272
rect 250444 369928 250496 369980
rect 337752 369928 337804 369980
rect 193128 369860 193180 369912
rect 337476 369860 337528 369912
rect 249064 367072 249116 367124
rect 337476 367072 337528 367124
rect 485044 364352 485096 364404
rect 580172 364352 580224 364404
rect 482284 351908 482336 351960
rect 580172 351908 580224 351960
rect 184848 349120 184900 349172
rect 337292 349120 337344 349172
rect 33048 347828 33100 347880
rect 37832 347828 37884 347880
rect 3056 345040 3108 345092
rect 32496 345040 32548 345092
rect 38108 339396 38160 339448
rect 131764 339396 131816 339448
rect 38292 339328 38344 339380
rect 153844 339328 153896 339380
rect 3424 339260 3476 339312
rect 132500 339260 132552 339312
rect 3516 339192 3568 339244
rect 136640 339192 136692 339244
rect 3608 339124 3660 339176
rect 140780 339124 140832 339176
rect 3792 339056 3844 339108
rect 155960 339056 156012 339108
rect 38844 338988 38896 339040
rect 193220 338988 193272 339040
rect 92296 338920 92348 338972
rect 580264 338920 580316 338972
rect 81348 338852 81400 338904
rect 580356 338852 580408 338904
rect 75828 338784 75880 338836
rect 580448 338784 580500 338836
rect 73068 338716 73120 338768
rect 580540 338716 580592 338768
rect 39764 338648 39816 338700
rect 126980 338648 127032 338700
rect 38568 338036 38620 338088
rect 337384 338036 337436 338088
rect 48964 337968 49016 338020
rect 368480 337968 368532 338020
rect 40500 337900 40552 337952
rect 356060 337900 356112 337952
rect 56508 337832 56560 337884
rect 236644 337832 236696 337884
rect 43444 337764 43496 337816
rect 394700 337764 394752 337816
rect 99288 337696 99340 337748
rect 226984 337696 227036 337748
rect 95148 337628 95200 337680
rect 225604 337628 225656 337680
rect 385684 337628 385736 337680
rect 387800 337628 387852 337680
rect 388444 337628 388496 337680
rect 390560 337628 390612 337680
rect 91008 337560 91060 337612
rect 239404 337560 239456 337612
rect 387064 337560 387116 337612
rect 389180 337560 389232 337612
rect 78588 337492 78640 337544
rect 239588 337492 239640 337544
rect 77208 337424 77260 337476
rect 239496 337424 239548 337476
rect 57888 337356 57940 337408
rect 221464 337356 221516 337408
rect 359464 337356 359516 337408
rect 378140 337356 378192 337408
rect 216588 337288 216640 337340
rect 382280 337288 382332 337340
rect 382924 337288 382976 337340
rect 390560 337288 390612 337340
rect 391296 337288 391348 337340
rect 397460 337288 397512 337340
rect 40408 337220 40460 337272
rect 59452 337220 59504 337272
rect 72976 337220 73028 337272
rect 239680 337220 239732 337272
rect 240048 337220 240100 337272
rect 398840 337220 398892 337272
rect 39396 337152 39448 337204
rect 59360 337152 59412 337204
rect 203524 337152 203576 337204
rect 371240 337152 371292 337204
rect 373264 337152 373316 337204
rect 445760 337152 445812 337204
rect 234528 337084 234580 337136
rect 396080 337084 396132 337136
rect 355324 337016 355376 337068
rect 375380 337016 375432 337068
rect 377404 337016 377456 337068
rect 391940 337016 391992 337068
rect 42064 336948 42116 337000
rect 361580 336948 361632 337000
rect 370504 336948 370556 337000
rect 437480 336948 437532 337000
rect 367744 336880 367796 336932
rect 434720 336880 434772 336932
rect 50344 336812 50396 336864
rect 369860 336812 369912 336864
rect 93584 336744 93636 336796
rect 100024 336744 100076 336796
rect 391204 336744 391256 336796
rect 393872 336744 393924 336796
rect 420184 336744 420236 336796
rect 422668 336744 422720 336796
rect 119988 336540 120040 336592
rect 178040 336540 178092 336592
rect 99288 336472 99340 336524
rect 171784 336472 171836 336524
rect 96528 336404 96580 336456
rect 173164 336404 173216 336456
rect 131028 336336 131080 336388
rect 213184 336336 213236 336388
rect 81256 336268 81308 336320
rect 177304 336268 177356 336320
rect 117228 336200 117280 336252
rect 214564 336200 214616 336252
rect 229744 336200 229796 336252
rect 385132 336200 385184 336252
rect 77208 336132 77260 336184
rect 242900 336132 242952 336184
rect 247684 336132 247736 336184
rect 369952 336132 370004 336184
rect 32404 336064 32456 336116
rect 143540 336064 143592 336116
rect 209688 336064 209740 336116
rect 400220 336064 400272 336116
rect 34428 335996 34480 336048
rect 382280 335996 382332 336048
rect 81072 334908 81124 334960
rect 200764 334908 200816 334960
rect 74908 334840 74960 334892
rect 195244 334840 195296 334892
rect 76288 334772 76340 334824
rect 243084 334772 243136 334824
rect 31392 334704 31444 334756
rect 386604 334704 386656 334756
rect 35716 334636 35768 334688
rect 396172 334636 396224 334688
rect 34336 334568 34388 334620
rect 407120 334568 407172 334620
rect 85304 333548 85356 333600
rect 162124 333548 162176 333600
rect 86408 333480 86460 333532
rect 169024 333480 169076 333532
rect 90640 333412 90692 333464
rect 220084 333412 220136 333464
rect 38660 333344 38712 333396
rect 189080 333344 189132 333396
rect 83556 333276 83608 333328
rect 244464 333276 244516 333328
rect 30288 333208 30340 333260
rect 360200 333208 360252 333260
rect 38660 324912 38712 324964
rect 67640 324912 67692 324964
rect 68836 324300 68888 324352
rect 580172 324300 580224 324352
rect 3424 318792 3476 318844
rect 156052 318792 156104 318844
rect 70308 311856 70360 311908
rect 580172 311856 580224 311908
rect 21456 311108 21508 311160
rect 150440 311108 150492 311160
rect 3424 304988 3476 305040
rect 158720 304988 158772 305040
rect 67548 298120 67600 298172
rect 580172 298120 580224 298172
rect 32864 297372 32916 297424
rect 387892 297372 387944 297424
rect 3424 292544 3476 292596
rect 157340 292544 157392 292596
rect 19984 290436 20036 290488
rect 146300 290436 146352 290488
rect 28264 282140 28316 282192
rect 139400 282140 139452 282192
rect 25504 280780 25556 280832
rect 149060 280780 149112 280832
rect 38752 277992 38804 278044
rect 241520 277992 241572 278044
rect 31668 275272 31720 275324
rect 364340 275272 364392 275324
rect 97908 273912 97960 273964
rect 232504 273912 232556 273964
rect 64696 271872 64748 271924
rect 579804 271872 579856 271924
rect 100024 271124 100076 271176
rect 230480 271124 230532 271176
rect 79968 269764 80020 269816
rect 244648 269764 244700 269816
rect 88156 268336 88208 268388
rect 167644 268336 167696 268388
rect 3056 266364 3108 266416
rect 160560 266364 160612 266416
rect 126888 265616 126940 265668
rect 222844 265616 222896 265668
rect 107568 264256 107620 264308
rect 262864 264256 262916 264308
rect 34244 264188 34296 264240
rect 380992 264188 381044 264240
rect 85488 262828 85540 262880
rect 196624 262828 196676 262880
rect 100024 261468 100076 261520
rect 527180 261468 527232 261520
rect 32496 260176 32548 260228
rect 154580 260176 154632 260228
rect 88156 260108 88208 260160
rect 258724 260108 258776 260160
rect 66168 258068 66220 258120
rect 580172 258068 580224 258120
rect 71688 257320 71740 257372
rect 482284 257320 482336 257372
rect 37004 255960 37056 256012
rect 92480 255960 92532 256012
rect 108764 255960 108816 256012
rect 333244 255960 333296 256012
rect 78496 254600 78548 254652
rect 244556 254600 244608 254652
rect 74356 254532 74408 254584
rect 245660 254532 245712 254584
rect 3424 253920 3476 253972
rect 163136 253920 163188 253972
rect 35808 253580 35860 253632
rect 135260 253580 135312 253632
rect 118608 253512 118660 253564
rect 220820 253512 220872 253564
rect 129648 253444 129700 253496
rect 243452 253444 243504 253496
rect 21364 253376 21416 253428
rect 148048 253376 148100 253428
rect 104716 253308 104768 253360
rect 327724 253308 327776 253360
rect 31484 253240 31536 253292
rect 367192 253240 367244 253292
rect 33968 253172 34020 253224
rect 409880 253172 409932 253224
rect 117964 252356 118016 252408
rect 201500 252356 201552 252408
rect 111616 252288 111668 252340
rect 211804 252288 211856 252340
rect 17224 252220 17276 252272
rect 135536 252220 135588 252272
rect 14464 252152 14516 252204
rect 153200 252152 153252 252204
rect 35440 252084 35492 252136
rect 113180 252084 113232 252136
rect 114468 252084 114520 252136
rect 266360 252084 266412 252136
rect 74448 252016 74500 252068
rect 243176 252016 243228 252068
rect 106096 251948 106148 252000
rect 334624 251948 334676 252000
rect 32680 251880 32732 251932
rect 383660 251880 383712 251932
rect 102048 251812 102100 251864
rect 480904 251812 480956 251864
rect 109500 251064 109552 251116
rect 193864 251064 193916 251116
rect 90732 250996 90784 251048
rect 189724 250996 189776 251048
rect 37096 250928 37148 250980
rect 142160 250928 142212 250980
rect 79416 250860 79468 250912
rect 185584 250860 185636 250912
rect 15844 250792 15896 250844
rect 132132 250792 132184 250844
rect 142068 250792 142120 250844
rect 242992 250792 243044 250844
rect 10324 250724 10376 250776
rect 142160 250724 142212 250776
rect 106188 250656 106240 250708
rect 240508 250656 240560 250708
rect 81900 250588 81952 250640
rect 255964 250588 256016 250640
rect 36912 250520 36964 250572
rect 100760 250520 100812 250572
rect 101956 250520 102008 250572
rect 330484 250520 330536 250572
rect 74448 250452 74500 250504
rect 483664 250452 483716 250504
rect 93216 249704 93268 249756
rect 182824 249704 182876 249756
rect 89444 249636 89496 249688
rect 180064 249636 180116 249688
rect 36728 249568 36780 249620
rect 122840 249568 122892 249620
rect 146208 249568 146260 249620
rect 239772 249568 239824 249620
rect 94504 249500 94556 249552
rect 191104 249500 191156 249552
rect 78220 249432 78272 249484
rect 178684 249432 178736 249484
rect 83188 249364 83240 249416
rect 186964 249364 187016 249416
rect 121368 249296 121420 249348
rect 240140 249296 240192 249348
rect 104808 249228 104860 249280
rect 240416 249228 240468 249280
rect 6184 249160 6236 249212
rect 130844 249160 130896 249212
rect 191104 249160 191156 249212
rect 359464 249160 359516 249212
rect 96988 249092 97040 249144
rect 479524 249092 479576 249144
rect 85672 249024 85724 249076
rect 545764 249024 545816 249076
rect 59268 247868 59320 247920
rect 187332 247868 187384 247920
rect 62028 247800 62080 247852
rect 241796 247800 241848 247852
rect 38108 247732 38160 247784
rect 261484 247732 261536 247784
rect 31576 247664 31628 247716
rect 358820 247664 358872 247716
rect 95700 246984 95752 247036
rect 207664 246984 207716 247036
rect 88248 246916 88300 246968
rect 204904 246916 204956 246968
rect 8208 246848 8260 246900
rect 128360 246848 128412 246900
rect 139308 246848 139360 246900
rect 240692 246848 240744 246900
rect 111708 246780 111760 246832
rect 240600 246780 240652 246832
rect 36820 246712 36872 246764
rect 107660 246712 107712 246764
rect 114560 246712 114612 246764
rect 282920 246712 282972 246764
rect 3700 246644 3752 246696
rect 152188 246644 152240 246696
rect 218152 246644 218204 246696
rect 412640 246644 412692 246696
rect 34060 246576 34112 246628
rect 372712 246576 372764 246628
rect 103244 246508 103296 246560
rect 477500 246508 477552 246560
rect 76932 246440 76984 246492
rect 486424 246440 486476 246492
rect 73160 246372 73212 246424
rect 485044 246372 485096 246424
rect 35072 246304 35124 246356
rect 70492 246304 70544 246356
rect 99472 246304 99524 246356
rect 542360 246304 542412 246356
rect 33784 246236 33836 246288
rect 143448 246236 143500 246288
rect 24768 246168 24820 246220
rect 129648 246168 129700 246220
rect 118332 246100 118384 246152
rect 218060 246100 218112 246152
rect 35164 245284 35216 245336
rect 134616 245284 134668 245336
rect 31024 245216 31076 245268
rect 138388 245216 138440 245268
rect 115848 245148 115900 245200
rect 234620 245148 234672 245200
rect 13084 245080 13136 245132
rect 145932 245080 145984 245132
rect 33784 245012 33836 245064
rect 168472 245012 168524 245064
rect 112076 244944 112128 244996
rect 299480 244944 299532 244996
rect 35256 244876 35308 244928
rect 172244 244876 172296 244928
rect 223672 244876 223724 244928
rect 420184 244876 420236 244928
rect 25504 244808 25556 244860
rect 164700 244808 164752 244860
rect 28264 244740 28316 244792
rect 176016 244740 176068 244792
rect 6184 244672 6236 244724
rect 179788 244672 179840 244724
rect 59360 244604 59412 244656
rect 265624 244604 265676 244656
rect 55588 244536 55640 244588
rect 262864 244536 262916 244588
rect 51816 244468 51868 244520
rect 261484 244468 261536 244520
rect 48044 244400 48096 244452
rect 258724 244400 258776 244452
rect 44272 244332 44324 244384
rect 255964 244332 256016 244384
rect 100760 244264 100812 244316
rect 579804 244264 579856 244316
rect 68100 244196 68152 244248
rect 68836 244196 68888 244248
rect 69388 244196 69440 244248
rect 70308 244196 70360 244248
rect 70676 244196 70728 244248
rect 71688 244196 71740 244248
rect 71872 244196 71924 244248
rect 73068 244196 73120 244248
rect 84476 244196 84528 244248
rect 85488 244196 85540 244248
rect 86960 244196 87012 244248
rect 88156 244196 88208 244248
rect 98276 244196 98328 244248
rect 100024 244196 100076 244248
rect 110788 244196 110840 244248
rect 111616 244196 111668 244248
rect 113272 244196 113324 244248
rect 114468 244196 114520 244248
rect 117044 244196 117096 244248
rect 117964 244196 118016 244248
rect 173164 244196 173216 244248
rect 7564 244128 7616 244180
rect 171048 244128 171100 244180
rect 171784 244128 171836 244180
rect 202328 244196 202380 244248
rect 203524 244196 203576 244248
rect 208676 244196 208728 244248
rect 209688 244196 209740 244248
rect 233700 244196 233752 244248
rect 234528 244196 234580 244248
rect 238760 244196 238812 244248
rect 240048 244196 240100 244248
rect 206100 244128 206152 244180
rect 213184 244128 213236 244180
rect 169024 244060 169076 244112
rect 222476 244060 222528 244112
rect 226984 244128 227036 244180
rect 236276 244128 236328 244180
rect 237472 244128 237524 244180
rect 373264 244128 373316 244180
rect 228732 244060 228784 244112
rect 229928 244060 229980 244112
rect 377404 244060 377456 244112
rect 162124 243992 162176 244044
rect 219900 243992 219952 244044
rect 224960 243992 225012 244044
rect 385684 243992 385736 244044
rect 153844 243924 153896 243976
rect 123300 243856 123352 243908
rect 176844 243856 176896 243908
rect 192300 243924 192352 243976
rect 193128 243924 193180 243976
rect 197360 243924 197412 243976
rect 198648 243924 198700 243976
rect 200764 243924 200816 243976
rect 213644 243924 213696 243976
rect 214932 243924 214984 243976
rect 380900 243924 380952 243976
rect 196072 243856 196124 243908
rect 207388 243856 207440 243908
rect 211160 243856 211212 243908
rect 122104 243788 122156 243840
rect 176752 243788 176804 243840
rect 214564 243788 214616 243840
rect 218704 243788 218756 243840
rect 63132 243720 63184 243772
rect 100760 243720 100812 243772
rect 120816 243720 120868 243772
rect 176660 243720 176712 243772
rect 177304 243720 177356 243772
rect 194876 243720 194928 243772
rect 195244 243720 195296 243772
rect 204904 243720 204956 243772
rect 376852 243856 376904 243908
rect 379612 243788 379664 243840
rect 379520 243720 379572 243772
rect 39672 243652 39724 243704
rect 124588 243652 124640 243704
rect 131764 243652 131816 243704
rect 198648 243652 198700 243704
rect 203616 243652 203668 243704
rect 374000 243652 374052 243704
rect 39856 243584 39908 243636
rect 125876 243584 125928 243636
rect 188528 243584 188580 243636
rect 363052 243584 363104 243636
rect 36636 243516 36688 243568
rect 132592 243516 132644 243568
rect 186044 243516 186096 243568
rect 362960 243516 363012 243568
rect 60648 243448 60700 243500
rect 115940 243448 115992 243500
rect 167644 243448 167696 243500
rect 201132 243448 201184 243500
rect 209872 243448 209924 243500
rect 225604 243448 225656 243500
rect 232228 243448 232280 243500
rect 61844 243380 61896 243432
rect 184664 243380 184716 243432
rect 199844 243380 199896 243432
rect 229744 243380 229796 243432
rect 46848 243312 46900 243364
rect 172428 243312 172480 243364
rect 183560 243312 183612 243364
rect 184848 243312 184900 243364
rect 212448 243312 212500 243364
rect 222844 243312 222896 243364
rect 226248 243312 226300 243364
rect 31760 243244 31812 243296
rect 162216 243244 162268 243296
rect 58072 243176 58124 243228
rect 187700 243176 187752 243228
rect 232504 243176 232556 243228
rect 234988 243176 235040 243228
rect 19984 243108 20036 243160
rect 167276 243108 167328 243160
rect 13084 243040 13136 243092
rect 174728 243040 174780 243092
rect 220084 243040 220136 243092
rect 227444 243040 227496 243092
rect 15844 242972 15896 243024
rect 178500 242972 178552 243024
rect 36544 242904 36596 242956
rect 40592 242904 40644 242956
rect 100760 242904 100812 242956
rect 102048 242904 102100 242956
rect 38568 242836 38620 242888
rect 39304 242836 39356 242888
rect 39856 242836 39908 242888
rect 91192 242836 91244 242888
rect 92388 242836 92440 242888
rect 240232 242836 240284 242888
rect 32772 242768 32824 242820
rect 70584 242768 70636 242820
rect 82728 242768 82780 242820
rect 243360 242768 243412 242820
rect 68928 242700 68980 242752
rect 243268 242700 243320 242752
rect 63408 242632 63460 242684
rect 240324 242632 240376 242684
rect 32956 242564 33008 242616
rect 337568 242564 337620 242616
rect 35532 242496 35584 242548
rect 376760 242496 376812 242548
rect 36452 242428 36504 242480
rect 385040 242428 385092 242480
rect 35348 242360 35400 242412
rect 420920 242360 420972 242412
rect 37188 242292 37240 242344
rect 440240 242292 440292 242344
rect 39212 242224 39264 242276
rect 443000 242224 443052 242276
rect 3424 242156 3476 242208
rect 31760 242156 31812 242208
rect 64788 242156 64840 242208
rect 244372 242156 244424 242208
rect 39028 242088 39080 242140
rect 88432 242088 88484 242140
rect 96344 242088 96396 242140
rect 244280 242088 244332 242140
rect 39948 242020 40000 242072
rect 98000 242020 98052 242072
rect 35624 241952 35676 242004
rect 82912 241952 82964 242004
rect 34152 241884 34204 241936
rect 69112 241884 69164 241936
rect 39120 241476 39172 241528
rect 39856 241476 39908 241528
rect 24124 241408 24176 241460
rect 173164 241408 173216 241460
rect 37832 241340 37884 241392
rect 43444 241340 43496 241392
rect 38292 241272 38344 241324
rect 48964 241272 49016 241324
rect 38568 241204 38620 241256
rect 42064 241204 42116 241256
rect 38844 241136 38896 241188
rect 37740 241068 37792 241120
rect 50344 241204 50396 241256
rect 57152 241247 57204 241256
rect 57152 241213 57161 241247
rect 57161 241213 57195 241247
rect 57195 241213 57204 241247
rect 57152 241204 57204 241213
rect 45928 241179 45980 241188
rect 43352 241111 43404 241120
rect 43352 241077 43361 241111
rect 43361 241077 43395 241111
rect 43395 241077 43404 241111
rect 43352 241068 43404 241077
rect 45928 241145 45937 241179
rect 45937 241145 45971 241179
rect 45971 241145 45980 241179
rect 45928 241136 45980 241145
rect 49608 241179 49660 241188
rect 49608 241145 49617 241179
rect 49617 241145 49651 241179
rect 49651 241145 49660 241179
rect 49608 241136 49660 241145
rect 50896 241179 50948 241188
rect 50896 241145 50905 241179
rect 50905 241145 50939 241179
rect 50939 241145 50948 241179
rect 50896 241136 50948 241145
rect 53472 241179 53524 241188
rect 53472 241145 53481 241179
rect 53481 241145 53515 241179
rect 53515 241145 53524 241179
rect 53472 241136 53524 241145
rect 54576 241179 54628 241188
rect 54576 241145 54585 241179
rect 54585 241145 54619 241179
rect 54619 241145 54628 241179
rect 54576 241136 54628 241145
rect 64972 241136 65024 241188
rect 115940 241179 115992 241188
rect 115940 241145 115949 241179
rect 115949 241145 115983 241179
rect 115983 241145 115992 241179
rect 115940 241136 115992 241145
rect 236644 241136 236696 241188
rect 241612 241136 241664 241188
rect 66352 241068 66404 241120
rect 83004 241111 83056 241120
rect 83004 241077 83013 241111
rect 83013 241077 83047 241111
rect 83047 241077 83056 241111
rect 83004 241068 83056 241077
rect 88064 241068 88116 241120
rect 241888 241068 241940 241120
rect 32404 241000 32456 241052
rect 165620 241000 165672 241052
rect 221464 241000 221516 241052
rect 241704 241000 241756 241052
rect 31024 240932 31076 240984
rect 169576 240932 169628 240984
rect 172428 240932 172480 240984
rect 21364 240864 21416 240916
rect 177028 240864 177080 240916
rect 38752 240796 38804 240848
rect 187700 240932 187752 240984
rect 580356 240932 580408 240984
rect 180892 240907 180944 240916
rect 180892 240873 180901 240907
rect 180901 240873 180935 240907
rect 180935 240873 180944 240907
rect 180892 240864 180944 240873
rect 182088 240907 182140 240916
rect 182088 240873 182097 240907
rect 182097 240873 182131 240907
rect 182131 240873 182140 240907
rect 182088 240864 182140 240873
rect 184664 240864 184716 240916
rect 580448 240864 580500 240916
rect 580264 240796 580316 240848
rect 38936 240728 38988 240780
rect 579804 240728 579856 240780
rect 14464 240660 14516 240712
rect 10324 240592 10376 240644
rect 273904 240524 273956 240576
rect 272524 240456 272576 240508
rect 269764 240388 269816 240440
rect 268384 240320 268436 240372
rect 280804 240252 280856 240304
rect 279424 240184 279476 240236
rect 276664 240116 276716 240168
rect 242808 234540 242860 234592
rect 391296 234540 391348 234592
rect 242808 223524 242860 223576
rect 367744 223524 367796 223576
rect 35808 217948 35860 218000
rect 38016 217948 38068 218000
rect 242808 217948 242860 218000
rect 388444 217948 388496 218000
rect 3332 215228 3384 215280
rect 25504 215228 25556 215280
rect 241980 212372 242032 212424
rect 243452 212372 243504 212424
rect 242532 208292 242584 208344
rect 427820 208292 427872 208344
rect 265624 206932 265676 206984
rect 579896 206932 579948 206984
rect 3424 202784 3476 202836
rect 19984 202784 20036 202836
rect 242440 202784 242492 202836
rect 387064 202784 387116 202836
rect 242348 197276 242400 197328
rect 424324 197276 424376 197328
rect 35348 195916 35400 195968
rect 38016 195916 38068 195968
rect 273904 193128 273956 193180
rect 580172 193128 580224 193180
rect 31392 191768 31444 191820
rect 38016 191768 38068 191820
rect 3424 188980 3476 189032
rect 32404 188980 32456 189032
rect 36452 187620 36504 187672
rect 37372 187620 37424 187672
rect 37832 186396 37884 186448
rect 40500 186396 40552 186448
rect 37096 186328 37148 186380
rect 37924 186328 37976 186380
rect 242808 186260 242860 186312
rect 386420 186260 386472 186312
rect 38384 183472 38436 183524
rect 39488 183472 39540 183524
rect 242808 180752 242860 180804
rect 417424 180752 417476 180804
rect 32680 177964 32732 178016
rect 38016 177964 38068 178016
rect 242808 175176 242860 175228
rect 415400 175176 415452 175228
rect 35440 173340 35492 173392
rect 38016 173340 38068 173392
rect 241888 169940 241940 169992
rect 244464 169940 244516 169992
rect 33968 169668 34020 169720
rect 38016 169668 38068 169720
rect 262864 166948 262916 167000
rect 580172 166948 580224 167000
rect 3240 164160 3292 164212
rect 33784 164160 33836 164212
rect 34336 161372 34388 161424
rect 38016 161372 38068 161424
rect 241888 159400 241940 159452
rect 243360 159400 243412 159452
rect 272524 153144 272576 153196
rect 579804 153144 579856 153196
rect 35532 151716 35584 151768
rect 38016 151716 38068 151768
rect 3424 150220 3476 150272
rect 7564 150220 7616 150272
rect 242808 148996 242860 149048
rect 405740 148996 405792 149048
rect 35716 147568 35768 147620
rect 38016 147568 38068 147620
rect 241888 143420 241940 143472
rect 244648 143420 244700 143472
rect 34060 139340 34112 139392
rect 38016 139340 38068 139392
rect 280804 139340 280856 139392
rect 580172 139340 580224 139392
rect 3240 137912 3292 137964
rect 31024 137912 31076 137964
rect 32864 131044 32916 131096
rect 38016 131044 38068 131096
rect 242256 128256 242308 128308
rect 393412 128256 393464 128308
rect 261484 126896 261536 126948
rect 580172 126896 580224 126948
rect 32772 125128 32824 125180
rect 38016 125128 38068 125180
rect 241980 122544 242032 122596
rect 245660 122544 245712 122596
rect 34152 121388 34204 121440
rect 37924 121388 37976 121440
rect 38200 117920 38252 117972
rect 39396 117920 39448 117972
rect 242808 117240 242860 117292
rect 254584 117240 254636 117292
rect 35624 113092 35676 113144
rect 38016 113092 38068 113144
rect 269764 113092 269816 113144
rect 580172 113092 580224 113144
rect 3424 111732 3476 111784
rect 35256 111732 35308 111784
rect 241888 111596 241940 111648
rect 243268 111596 243320 111648
rect 34428 108944 34480 108996
rect 37648 108944 37700 108996
rect 241888 107516 241940 107568
rect 244556 107516 244608 107568
rect 279424 100648 279476 100700
rect 580172 100648 580224 100700
rect 3424 97928 3476 97980
rect 13084 97928 13136 97980
rect 242808 95956 242860 96008
rect 250444 95956 250496 96008
rect 34244 95140 34296 95192
rect 38016 95140 38068 95192
rect 31484 90992 31536 91044
rect 38016 90992 38068 91044
rect 258724 86912 258776 86964
rect 580172 86912 580224 86964
rect 3148 85484 3200 85536
rect 24124 85484 24176 85536
rect 242256 79976 242308 80028
rect 249064 79976 249116 80028
rect 30288 76916 30340 76968
rect 38016 76916 38068 76968
rect 241520 74468 241572 74520
rect 243176 74468 243228 74520
rect 268384 73108 268436 73160
rect 579988 73108 580040 73160
rect 3424 71680 3476 71732
rect 28264 71680 28316 71732
rect 31668 68960 31720 69012
rect 38016 68960 38068 69012
rect 242808 64812 242860 64864
rect 356152 64812 356204 64864
rect 31576 60664 31628 60716
rect 38016 60664 38068 60716
rect 3056 59304 3108 59356
rect 15844 59304 15896 59356
rect 241520 58896 241572 58948
rect 244372 58896 244424 58948
rect 35072 56516 35124 56568
rect 38016 56516 38068 56568
rect 241980 53728 242032 53780
rect 357440 53728 357492 53780
rect 32956 46860 33008 46912
rect 38016 46860 38068 46912
rect 255964 46860 256016 46912
rect 580172 46860 580224 46912
rect 3424 45500 3476 45552
rect 21364 45500 21416 45552
rect 33048 42712 33100 42764
rect 38016 42712 38068 42764
rect 36544 39312 36596 39364
rect 580264 39312 580316 39364
rect 220176 39040 220228 39092
rect 355324 39040 355376 39092
rect 232964 38972 233016 39024
rect 392584 38972 392636 39024
rect 200212 38904 200264 38956
rect 367100 38904 367152 38956
rect 223028 38836 223080 38888
rect 397552 38836 397604 38888
rect 225880 38768 225932 38820
rect 402980 38768 403032 38820
rect 230112 38700 230164 38752
rect 430580 38700 430632 38752
rect 38476 38632 38528 38684
rect 215852 38632 215904 38684
rect 231584 38632 231636 38684
rect 433340 38632 433392 38684
rect 39304 38564 39356 38616
rect 40684 38564 40736 38616
rect 195888 38564 195940 38616
rect 237288 38564 237340 38616
rect 244280 38564 244332 38616
rect 37096 38496 37148 38548
rect 213000 38496 213052 38548
rect 224408 38496 224460 38548
rect 239588 38496 239640 38548
rect 40408 38428 40460 38480
rect 204444 38428 204496 38480
rect 227260 38428 227312 38480
rect 240140 38428 240192 38480
rect 39488 38360 39540 38412
rect 197360 38360 197412 38412
rect 228732 38360 228784 38412
rect 240232 38360 240284 38412
rect 207296 38292 207348 38344
rect 365720 38292 365772 38344
rect 60004 38224 60056 38276
rect 69112 38224 69164 38276
rect 90364 38224 90416 38276
rect 147496 38224 147548 38276
rect 151084 38224 151136 38276
rect 160284 38224 160336 38276
rect 234436 38224 234488 38276
rect 391204 38224 391256 38276
rect 66904 38156 66956 38208
rect 79140 38156 79192 38208
rect 61384 38088 61436 38140
rect 74816 38088 74868 38140
rect 79324 38088 79376 38140
rect 91928 38088 91980 38140
rect 37096 38020 37148 38072
rect 83372 38020 83424 38072
rect 39948 37952 40000 38004
rect 87696 37952 87748 38004
rect 46848 37884 46900 37936
rect 96160 37884 96212 37936
rect 100024 37884 100076 37936
rect 156052 38156 156104 38208
rect 160744 38156 160796 38208
rect 165988 38156 166040 38208
rect 201592 38156 201644 38208
rect 247684 38156 247736 38208
rect 108304 38088 108356 38140
rect 168840 38088 168892 38140
rect 169024 38088 169076 38140
rect 178868 38088 178920 38140
rect 208768 38088 208820 38140
rect 251824 38088 251876 38140
rect 104164 38020 104216 38072
rect 164608 38020 164660 38072
rect 164884 38020 164936 38072
rect 170312 38020 170364 38072
rect 175924 38020 175976 38072
rect 188804 38020 188856 38072
rect 221556 38020 221608 38072
rect 239496 38020 239548 38072
rect 104900 37952 104952 38004
rect 106188 37952 106240 38004
rect 106280 37952 106332 38004
rect 107568 37952 107620 38004
rect 115204 37952 115256 38004
rect 177396 37952 177448 38004
rect 178684 37952 178736 38004
rect 190276 37952 190328 38004
rect 205916 37952 205968 38004
rect 375472 37952 375524 38004
rect 122104 37884 122156 37936
rect 185952 37884 186004 37936
rect 217324 37884 217376 37936
rect 382924 37884 382976 37936
rect 51724 37816 51776 37868
rect 53472 37816 53524 37868
rect 57980 37816 58032 37868
rect 59176 37816 59228 37868
rect 60740 37816 60792 37868
rect 62028 37816 62080 37868
rect 149060 37816 149112 37868
rect 150348 37816 150400 37868
rect 172612 37816 172664 37868
rect 174544 37816 174596 37868
rect 203064 37816 203116 37868
rect 371884 37816 371936 37868
rect 211620 37748 211672 37800
rect 371332 37748 371384 37800
rect 55864 37680 55916 37732
rect 63408 37680 63460 37732
rect 69664 37680 69716 37732
rect 70584 37680 70636 37732
rect 113824 37680 113876 37732
rect 114744 37680 114796 37732
rect 147680 37680 147732 37732
rect 148876 37680 148928 37732
rect 174544 37680 174596 37732
rect 180248 37680 180300 37732
rect 214472 37680 214524 37732
rect 239680 37680 239732 37732
rect 218704 37612 218756 37664
rect 239404 37612 239456 37664
rect 238668 37544 238720 37596
rect 242992 37544 243044 37596
rect 48964 37476 49016 37528
rect 52000 37476 52052 37528
rect 146944 37408 146996 37460
rect 151728 37408 151780 37460
rect 54484 37272 54536 37324
rect 57704 37272 57756 37324
rect 177304 37272 177356 37324
rect 181720 37272 181772 37324
rect 19984 37136 20036 37188
rect 54852 37136 54904 37188
rect 75184 37136 75236 37188
rect 99012 37136 99064 37188
rect 8208 37068 8260 37120
rect 49148 37068 49200 37120
rect 73804 37068 73856 37120
rect 103336 37068 103388 37120
rect 32404 37000 32456 37052
rect 76288 37000 76340 37052
rect 82084 37000 82136 37052
rect 111892 37000 111944 37052
rect 34428 36932 34480 36984
rect 80520 36932 80572 36984
rect 83464 36932 83516 36984
rect 130384 36932 130436 36984
rect 15844 36864 15896 36916
rect 43352 36864 43404 36916
rect 43444 36864 43496 36916
rect 90548 36864 90600 36916
rect 95884 36864 95936 36916
rect 113272 36864 113324 36916
rect 38568 36796 38620 36848
rect 86224 36796 86276 36848
rect 91744 36796 91796 36848
rect 116124 36796 116176 36848
rect 4068 36728 4120 36780
rect 44916 36728 44968 36780
rect 53748 36728 53800 36780
rect 104716 36728 104768 36780
rect 17868 36660 17920 36712
rect 60556 36660 60608 36712
rect 68284 36660 68336 36712
rect 118976 36660 119028 36712
rect 22008 36592 22060 36644
rect 66260 36592 66312 36644
rect 71044 36592 71096 36644
rect 123300 36592 123352 36644
rect 123484 36592 123536 36644
rect 176016 36592 176068 36644
rect 2044 36524 2096 36576
rect 40684 36524 40736 36576
rect 57888 36524 57940 36576
rect 109040 36524 109092 36576
rect 119988 36524 120040 36576
rect 184572 36524 184624 36576
rect 87604 35912 87656 35964
rect 94780 35912 94832 35964
rect 126244 35912 126296 35964
rect 134708 35912 134760 35964
rect 25504 35504 25556 35556
rect 60740 35504 60792 35556
rect 35808 35436 35860 35488
rect 81992 35436 82044 35488
rect 28908 35368 28960 35420
rect 73436 35368 73488 35420
rect 77944 35368 77996 35420
rect 126152 35368 126204 35420
rect 24124 35300 24176 35352
rect 50620 35300 50672 35352
rect 50988 35300 51040 35352
rect 99380 35300 99432 35352
rect 31668 35232 31720 35284
rect 77668 35232 77720 35284
rect 86224 35232 86276 35284
rect 138940 35232 138992 35284
rect 13728 35164 13780 35216
rect 55220 35164 55272 35216
rect 64788 35164 64840 35216
rect 117596 35164 117648 35216
rect 117964 34484 118016 34536
rect 121828 34484 121880 34536
rect 267004 33056 267056 33108
rect 580172 33056 580224 33108
rect 2780 32784 2832 32836
rect 6184 32784 6236 32836
rect 6276 32376 6328 32428
rect 46296 32376 46348 32428
rect 111708 29588 111760 29640
rect 172612 29588 172664 29640
rect 3424 20612 3476 20664
rect 14464 20612 14516 20664
rect 276664 20612 276716 20664
rect 580172 20612 580224 20664
rect 88248 8916 88300 8968
rect 132500 8916 132552 8968
rect 24768 7556 24820 7608
rect 67640 7556 67692 7608
rect 95332 7556 95384 7608
rect 153200 7556 153252 7608
rect 3424 6808 3476 6860
rect 10324 6808 10376 6860
rect 85212 6604 85264 6656
rect 136640 6604 136692 6656
rect 61660 6536 61712 6588
rect 110420 6536 110472 6588
rect 115296 6536 115348 6588
rect 169024 6536 169076 6588
rect 108120 6468 108172 6520
rect 164884 6468 164936 6520
rect 104532 6400 104584 6452
rect 160744 6400 160796 6452
rect 51356 6332 51408 6384
rect 100760 6332 100812 6384
rect 101036 6332 101088 6384
rect 161480 6332 161532 6384
rect 47860 6264 47912 6316
rect 96620 6264 96672 6316
rect 97448 6264 97500 6316
rect 157340 6264 157392 6316
rect 54944 6196 54996 6248
rect 104900 6196 104952 6248
rect 118792 6196 118844 6248
rect 182180 6196 182232 6248
rect 62028 6128 62080 6180
rect 113824 6128 113876 6180
rect 122288 6128 122340 6180
rect 186320 6128 186372 6180
rect 76196 5448 76248 5500
rect 131120 5448 131172 5500
rect 72608 5380 72660 5432
rect 126980 5380 127032 5432
rect 70308 5312 70360 5364
rect 124220 5312 124272 5364
rect 79692 5244 79744 5296
rect 135260 5244 135312 5296
rect 83280 5176 83332 5228
rect 139400 5176 139452 5228
rect 86868 5108 86920 5160
rect 143540 5108 143592 5160
rect 90456 5040 90508 5092
rect 147680 5040 147732 5092
rect 29000 4972 29052 5024
rect 71780 4972 71832 5024
rect 87972 4972 88024 5024
rect 144920 4972 144972 5024
rect 40684 4904 40736 4956
rect 88340 4904 88392 4956
rect 102232 4904 102284 4956
rect 162860 4904 162912 4956
rect 37188 4836 37240 4888
rect 84200 4836 84252 4888
rect 95148 4836 95200 4888
rect 154580 4836 154632 4888
rect 9956 4768 10008 4820
rect 48964 4768 49016 4820
rect 56048 4768 56100 4820
rect 106280 4768 106332 4820
rect 109316 4768 109368 4820
rect 171140 4768 171192 4820
rect 73804 4700 73856 4752
rect 128360 4700 128412 4752
rect 66720 4632 66772 4684
rect 120080 4632 120132 4684
rect 43076 4088 43128 4140
rect 79324 4088 79376 4140
rect 103336 4088 103388 4140
rect 104164 4088 104216 4140
rect 123484 4088 123536 4140
rect 175924 4088 175976 4140
rect 19432 4020 19484 4072
rect 54484 4020 54536 4072
rect 24216 3952 24268 4004
rect 60004 3952 60056 4004
rect 63224 3952 63276 4004
rect 91744 4020 91796 4072
rect 92756 4020 92808 4072
rect 146944 4020 146996 4072
rect 67916 3952 67968 4004
rect 117964 3952 118016 4004
rect 124680 3952 124732 4004
rect 178684 3952 178736 4004
rect 11152 3884 11204 3936
rect 51724 3884 51776 3936
rect 52552 3884 52604 3936
rect 73712 3884 73764 3936
rect 85672 3884 85724 3936
rect 142160 3884 142212 3936
rect 14740 3816 14792 3868
rect 55864 3816 55916 3868
rect 59636 3816 59688 3868
rect 81992 3816 82044 3868
rect 82084 3816 82136 3868
rect 6460 3748 6512 3800
rect 46940 3748 46992 3800
rect 48964 3748 49016 3800
rect 84476 3816 84528 3868
rect 140780 3816 140832 3868
rect 86224 3748 86276 3800
rect 91560 3748 91612 3800
rect 149060 3748 149112 3800
rect 15936 3680 15988 3732
rect 57980 3680 58032 3732
rect 60832 3680 60884 3732
rect 95884 3680 95936 3732
rect 117596 3680 117648 3732
rect 30104 3612 30156 3664
rect 32404 3612 32456 3664
rect 45468 3612 45520 3664
rect 87604 3612 87656 3664
rect 114008 3612 114060 3664
rect 115204 3612 115256 3664
rect 121092 3612 121144 3664
rect 122104 3612 122156 3664
rect 174544 3680 174596 3732
rect 177304 3612 177356 3664
rect 1676 3544 1728 3596
rect 10324 3544 10376 3596
rect 12348 3544 12400 3596
rect 19984 3544 20036 3596
rect 25320 3544 25372 3596
rect 69664 3544 69716 3596
rect 75000 3544 75052 3596
rect 83464 3544 83516 3596
rect 98644 3544 98696 3596
rect 158720 3544 158772 3596
rect 193128 3544 193180 3596
rect 582196 3544 582248 3596
rect 5264 3476 5316 3528
rect 6276 3476 6328 3528
rect 7656 3476 7708 3528
rect 8208 3476 8260 3528
rect 17040 3476 17092 3528
rect 17868 3476 17920 3528
rect 23020 3476 23072 3528
rect 24768 3476 24820 3528
rect 2872 3408 2924 3460
rect 15844 3408 15896 3460
rect 20628 3408 20680 3460
rect 64880 3476 64932 3528
rect 65524 3476 65576 3528
rect 68284 3476 68336 3528
rect 69112 3476 69164 3528
rect 71044 3476 71096 3528
rect 77392 3476 77444 3528
rect 88248 3476 88300 3528
rect 89168 3476 89220 3528
rect 90364 3476 90416 3528
rect 93952 3476 94004 3528
rect 95332 3476 95384 3528
rect 106924 3476 106976 3528
rect 108304 3476 108356 3528
rect 110512 3476 110564 3528
rect 172520 3476 172572 3528
rect 194508 3476 194560 3528
rect 583392 3476 583444 3528
rect 27712 3408 27764 3460
rect 28908 3408 28960 3460
rect 33600 3408 33652 3460
rect 34428 3408 34480 3460
rect 34796 3408 34848 3460
rect 35808 3408 35860 3460
rect 35992 3408 36044 3460
rect 37096 3408 37148 3460
rect 41880 3408 41932 3460
rect 43444 3408 43496 3460
rect 44272 3408 44324 3460
rect 92480 3408 92532 3460
rect 105728 3408 105780 3460
rect 167000 3408 167052 3460
rect 191748 3408 191800 3460
rect 581000 3408 581052 3460
rect 572 3340 624 3392
rect 2044 3340 2096 3392
rect 8760 3340 8812 3392
rect 24124 3340 24176 3392
rect 32404 3340 32456 3392
rect 66904 3340 66956 3392
rect 71504 3340 71556 3392
rect 77944 3340 77996 3392
rect 80888 3340 80940 3392
rect 85212 3340 85264 3392
rect 99840 3340 99892 3392
rect 151084 3340 151136 3392
rect 28908 3272 28960 3324
rect 50160 3272 50212 3324
rect 50988 3272 51040 3324
rect 57244 3272 57296 3324
rect 57888 3272 57940 3324
rect 58440 3272 58492 3324
rect 61660 3272 61712 3324
rect 64328 3272 64380 3324
rect 64788 3272 64840 3324
rect 75184 3272 75236 3324
rect 78588 3272 78640 3324
rect 126244 3272 126296 3324
rect 61384 3204 61436 3256
rect 112812 3204 112864 3256
rect 123392 3204 123444 3256
rect 96252 3136 96304 3188
rect 100024 3136 100076 3188
rect 116400 3136 116452 3188
rect 18236 2864 18288 2916
rect 25504 2864 25556 2916
rect 26516 2796 26568 2848
rect 29000 2796 29052 2848
<< metal2 >>
rect 8086 703520 8198 704960
rect 24278 703520 24390 704960
rect 40470 703520 40582 704960
rect 56754 703520 56866 704960
rect 72946 703520 73058 704960
rect 89138 703520 89250 704960
rect 105422 703520 105534 704960
rect 121614 703520 121726 704960
rect 137806 703520 137918 704960
rect 154090 703520 154202 704960
rect 170282 703520 170394 704960
rect 186474 703520 186586 704960
rect 202758 703520 202870 704960
rect 218072 703582 218836 703610
rect 8128 702434 8156 703520
rect 8128 702406 8248 702434
rect 2778 684312 2834 684321
rect 2778 684247 2834 684256
rect 2792 683670 2820 684247
rect 2780 683664 2832 683670
rect 2780 683606 2832 683612
rect 6184 683664 6236 683670
rect 6184 683606 6236 683612
rect 3422 671256 3478 671265
rect 3422 671191 3478 671200
rect 3330 606112 3386 606121
rect 3330 606047 3386 606056
rect 3344 605878 3372 606047
rect 3332 605872 3384 605878
rect 3332 605814 3384 605820
rect 3330 580000 3386 580009
rect 3330 579935 3386 579944
rect 3344 579698 3372 579935
rect 3332 579692 3384 579698
rect 3332 579634 3384 579640
rect 3330 553888 3386 553897
rect 3330 553823 3386 553832
rect 3344 553450 3372 553823
rect 3332 553444 3384 553450
rect 3332 553386 3384 553392
rect 3330 527912 3386 527921
rect 3330 527847 3386 527856
rect 3344 527202 3372 527847
rect 3332 527196 3384 527202
rect 3332 527138 3384 527144
rect 3330 514856 3386 514865
rect 3330 514791 3332 514800
rect 3384 514791 3386 514800
rect 3332 514762 3384 514768
rect 2870 501800 2926 501809
rect 2870 501735 2926 501744
rect 2884 501022 2912 501735
rect 2872 501016 2924 501022
rect 2872 500958 2924 500964
rect 3330 475688 3386 475697
rect 3330 475623 3386 475632
rect 3344 474774 3372 475623
rect 3332 474768 3384 474774
rect 3332 474710 3384 474716
rect 3330 462632 3386 462641
rect 3330 462567 3386 462576
rect 3344 462398 3372 462567
rect 3332 462392 3384 462398
rect 3332 462334 3384 462340
rect 3330 449576 3386 449585
rect 3330 449511 3386 449520
rect 3344 448594 3372 449511
rect 3332 448588 3384 448594
rect 3332 448530 3384 448536
rect 3146 423600 3202 423609
rect 3146 423535 3202 423544
rect 3160 422346 3188 423535
rect 3148 422340 3200 422346
rect 3148 422282 3200 422288
rect 3332 397520 3384 397526
rect 3330 397488 3332 397497
rect 3384 397488 3386 397497
rect 3330 397423 3386 397432
rect 3330 371376 3386 371385
rect 3330 371311 3386 371320
rect 3344 371278 3372 371311
rect 3332 371272 3384 371278
rect 3332 371214 3384 371220
rect 3054 345400 3110 345409
rect 3054 345335 3110 345344
rect 3068 345098 3096 345335
rect 3056 345092 3108 345098
rect 3056 345034 3108 345040
rect 3436 339318 3464 671191
rect 3514 658200 3570 658209
rect 3514 658135 3570 658144
rect 3528 656946 3556 658135
rect 3516 656940 3568 656946
rect 3516 656882 3568 656888
rect 3516 632120 3568 632126
rect 3514 632088 3516 632097
rect 3568 632088 3570 632097
rect 3514 632023 3570 632032
rect 3514 619168 3570 619177
rect 3514 619103 3570 619112
rect 3424 339312 3476 339318
rect 3424 339254 3476 339260
rect 3528 339250 3556 619103
rect 3606 566944 3662 566953
rect 3606 566879 3662 566888
rect 3516 339244 3568 339250
rect 3516 339186 3568 339192
rect 3620 339182 3648 566879
rect 3698 410544 3754 410553
rect 3698 410479 3754 410488
rect 3608 339176 3660 339182
rect 3608 339118 3660 339124
rect 3422 319288 3478 319297
rect 3422 319223 3478 319232
rect 3436 318850 3464 319223
rect 3424 318844 3476 318850
rect 3424 318786 3476 318792
rect 3422 306232 3478 306241
rect 3422 306167 3478 306176
rect 3436 305046 3464 306167
rect 3424 305040 3476 305046
rect 3424 304982 3476 304988
rect 3422 293176 3478 293185
rect 3422 293111 3478 293120
rect 3436 292602 3464 293111
rect 3424 292596 3476 292602
rect 3424 292538 3476 292544
rect 3054 267200 3110 267209
rect 3054 267135 3110 267144
rect 3068 266422 3096 267135
rect 3056 266416 3108 266422
rect 3056 266358 3108 266364
rect 3422 254144 3478 254153
rect 3422 254079 3478 254088
rect 3436 253978 3464 254079
rect 3424 253972 3476 253978
rect 3424 253914 3476 253920
rect 3712 246702 3740 410479
rect 3790 358456 3846 358465
rect 3790 358391 3846 358400
rect 3804 339114 3832 358391
rect 3792 339108 3844 339114
rect 3792 339050 3844 339056
rect 6196 249218 6224 683606
rect 6184 249212 6236 249218
rect 6184 249154 6236 249160
rect 8220 246906 8248 702406
rect 24320 699718 24348 703520
rect 39856 700324 39908 700330
rect 39856 700266 39908 700272
rect 24308 699712 24360 699718
rect 24308 699654 24360 699660
rect 24768 699712 24820 699718
rect 24768 699654 24820 699660
rect 39764 699712 39816 699718
rect 39764 699654 39816 699660
rect 15844 656940 15896 656946
rect 15844 656882 15896 656888
rect 10324 527196 10376 527202
rect 10324 527138 10376 527144
rect 10336 250782 10364 527138
rect 13084 474768 13136 474774
rect 13084 474710 13136 474716
rect 10324 250776 10376 250782
rect 10324 250718 10376 250724
rect 8208 246900 8260 246906
rect 8208 246842 8260 246848
rect 3700 246696 3752 246702
rect 3700 246638 3752 246644
rect 13096 245138 13124 474710
rect 14464 371272 14516 371278
rect 14464 371214 14516 371220
rect 14476 252210 14504 371214
rect 14464 252204 14516 252210
rect 14464 252146 14516 252152
rect 15856 250850 15884 656882
rect 17224 605872 17276 605878
rect 17224 605814 17276 605820
rect 17236 252278 17264 605814
rect 21364 462392 21416 462398
rect 21364 462334 21416 462340
rect 19984 448588 20036 448594
rect 19984 448530 20036 448536
rect 19996 290494 20024 448530
rect 19984 290488 20036 290494
rect 19984 290430 20036 290436
rect 21376 253434 21404 462334
rect 21456 397520 21508 397526
rect 21456 397462 21508 397468
rect 21468 311166 21496 397462
rect 21456 311160 21508 311166
rect 21456 311102 21508 311108
rect 21364 253428 21416 253434
rect 21364 253370 21416 253376
rect 17224 252272 17276 252278
rect 17224 252214 17276 252220
rect 15844 250844 15896 250850
rect 15844 250786 15896 250792
rect 24780 246226 24808 699654
rect 35164 632120 35216 632126
rect 35164 632062 35216 632068
rect 31024 579692 31076 579698
rect 31024 579634 31076 579640
rect 28264 553444 28316 553450
rect 28264 553386 28316 553392
rect 25504 422340 25556 422346
rect 25504 422282 25556 422288
rect 25516 280838 25544 422282
rect 28276 282198 28304 553386
rect 30288 333260 30340 333266
rect 30288 333202 30340 333208
rect 28264 282192 28316 282198
rect 28264 282134 28316 282140
rect 25504 280832 25556 280838
rect 25504 280774 25556 280780
rect 24768 246220 24820 246226
rect 24768 246162 24820 246168
rect 13084 245132 13136 245138
rect 13084 245074 13136 245080
rect 25504 244860 25556 244866
rect 25504 244802 25556 244808
rect 6184 244724 6236 244730
rect 6184 244666 6236 244672
rect 3424 242208 3476 242214
rect 3424 242150 3476 242156
rect 3436 241097 3464 242150
rect 3422 241088 3478 241097
rect 3422 241023 3478 241032
rect 3332 215280 3384 215286
rect 3332 215222 3384 215228
rect 3344 214985 3372 215222
rect 3330 214976 3386 214985
rect 3330 214911 3386 214920
rect 3424 202836 3476 202842
rect 3424 202778 3476 202784
rect 3436 201929 3464 202778
rect 3422 201920 3478 201929
rect 3422 201855 3478 201864
rect 3424 189032 3476 189038
rect 3424 188974 3476 188980
rect 3436 188873 3464 188974
rect 3422 188864 3478 188873
rect 3422 188799 3478 188808
rect 3240 164212 3292 164218
rect 3240 164154 3292 164160
rect 3252 162897 3280 164154
rect 3238 162888 3294 162897
rect 3238 162823 3294 162832
rect 3424 150272 3476 150278
rect 3424 150214 3476 150220
rect 3436 149841 3464 150214
rect 3422 149832 3478 149841
rect 3422 149767 3478 149776
rect 3240 137964 3292 137970
rect 3240 137906 3292 137912
rect 3252 136785 3280 137906
rect 3238 136776 3294 136785
rect 3238 136711 3294 136720
rect 3424 111784 3476 111790
rect 3424 111726 3476 111732
rect 3436 110673 3464 111726
rect 3422 110664 3478 110673
rect 3422 110599 3478 110608
rect 3424 97980 3476 97986
rect 3424 97922 3476 97928
rect 3436 97617 3464 97922
rect 3422 97608 3478 97617
rect 3422 97543 3478 97552
rect 3148 85536 3200 85542
rect 3148 85478 3200 85484
rect 3160 84697 3188 85478
rect 3146 84688 3202 84697
rect 3146 84623 3202 84632
rect 3424 71732 3476 71738
rect 3424 71674 3476 71680
rect 3436 71641 3464 71674
rect 3422 71632 3478 71641
rect 3422 71567 3478 71576
rect 3056 59356 3108 59362
rect 3056 59298 3108 59304
rect 3068 58585 3096 59298
rect 3054 58576 3110 58585
rect 3054 58511 3110 58520
rect 3424 45552 3476 45558
rect 3422 45520 3424 45529
rect 3476 45520 3478 45529
rect 3422 45455 3478 45464
rect 4068 36780 4120 36786
rect 4068 36722 4120 36728
rect 2044 36576 2096 36582
rect 2044 36518 2096 36524
rect 1676 3596 1728 3602
rect 1676 3538 1728 3544
rect 572 3392 624 3398
rect 572 3334 624 3340
rect 584 480 612 3334
rect 1688 480 1716 3538
rect 2056 3398 2084 36518
rect 2780 32836 2832 32842
rect 2780 32778 2832 32784
rect 2792 32473 2820 32778
rect 2778 32464 2834 32473
rect 2778 32399 2834 32408
rect 3424 20664 3476 20670
rect 3424 20606 3476 20612
rect 3436 19417 3464 20606
rect 3422 19408 3478 19417
rect 3422 19343 3478 19352
rect 3424 6860 3476 6866
rect 3424 6802 3476 6808
rect 3436 6497 3464 6802
rect 3422 6488 3478 6497
rect 3422 6423 3478 6432
rect 2872 3460 2924 3466
rect 2872 3402 2924 3408
rect 2044 3392 2096 3398
rect 2044 3334 2096 3340
rect 2884 480 2912 3402
rect 4080 480 4108 36722
rect 6196 32842 6224 244666
rect 7564 244180 7616 244186
rect 7564 244122 7616 244128
rect 7576 150278 7604 244122
rect 19984 243160 20036 243166
rect 19984 243102 20036 243108
rect 13084 243092 13136 243098
rect 13084 243034 13136 243040
rect 10324 240644 10376 240650
rect 10324 240586 10376 240592
rect 7564 150272 7616 150278
rect 7564 150214 7616 150220
rect 8208 37120 8260 37126
rect 8208 37062 8260 37068
rect 6184 32836 6236 32842
rect 6184 32778 6236 32784
rect 6276 32428 6328 32434
rect 6276 32370 6328 32376
rect 6288 3534 6316 32370
rect 6460 3800 6512 3806
rect 6460 3742 6512 3748
rect 5264 3528 5316 3534
rect 5264 3470 5316 3476
rect 6276 3528 6328 3534
rect 6276 3470 6328 3476
rect 5276 480 5304 3470
rect 6472 480 6500 3742
rect 8220 3534 8248 37062
rect 10336 6866 10364 240586
rect 13096 97986 13124 243034
rect 15844 243024 15896 243030
rect 15844 242966 15896 242972
rect 14464 240712 14516 240718
rect 14464 240654 14516 240660
rect 13084 97980 13136 97986
rect 13084 97922 13136 97928
rect 13728 35216 13780 35222
rect 13728 35158 13780 35164
rect 13740 6914 13768 35158
rect 14476 20670 14504 240654
rect 15856 59362 15884 242966
rect 19996 202842 20024 243102
rect 24124 241460 24176 241466
rect 24124 241402 24176 241408
rect 21364 240916 21416 240922
rect 21364 240858 21416 240864
rect 19984 202836 20036 202842
rect 19984 202778 20036 202784
rect 15844 59356 15896 59362
rect 15844 59298 15896 59304
rect 21376 45558 21404 240858
rect 24136 85542 24164 241402
rect 25516 215286 25544 244802
rect 28264 244792 28316 244798
rect 28264 244734 28316 244740
rect 25504 215280 25556 215286
rect 25504 215222 25556 215228
rect 24124 85536 24176 85542
rect 24124 85478 24176 85484
rect 28276 71738 28304 244734
rect 30300 76974 30328 333202
rect 31036 245274 31064 579634
rect 32404 514820 32456 514826
rect 32404 514762 32456 514768
rect 32416 336122 32444 514762
rect 33784 501016 33836 501022
rect 33784 500958 33836 500964
rect 33048 347880 33100 347886
rect 33048 347822 33100 347828
rect 32496 345092 32548 345098
rect 32496 345034 32548 345040
rect 32404 336116 32456 336122
rect 32404 336058 32456 336064
rect 31392 334756 31444 334762
rect 31392 334698 31444 334704
rect 31024 245268 31076 245274
rect 31024 245210 31076 245216
rect 31024 240984 31076 240990
rect 31024 240926 31076 240932
rect 31036 137970 31064 240926
rect 31404 191826 31432 334698
rect 31668 275324 31720 275330
rect 31668 275266 31720 275272
rect 31484 253292 31536 253298
rect 31484 253234 31536 253240
rect 31392 191820 31444 191826
rect 31392 191762 31444 191768
rect 31024 137964 31076 137970
rect 31024 137906 31076 137912
rect 31496 91050 31524 253234
rect 31576 247716 31628 247722
rect 31576 247658 31628 247664
rect 31484 91044 31536 91050
rect 31484 90986 31536 90992
rect 30288 76968 30340 76974
rect 30288 76910 30340 76916
rect 28264 71732 28316 71738
rect 28264 71674 28316 71680
rect 31588 60722 31616 247658
rect 31680 69018 31708 275266
rect 32508 260234 32536 345034
rect 32864 297424 32916 297430
rect 32864 297366 32916 297372
rect 32496 260228 32548 260234
rect 32496 260170 32548 260176
rect 32680 251932 32732 251938
rect 32680 251874 32732 251880
rect 31760 243296 31812 243302
rect 31760 243238 31812 243244
rect 31772 242214 31800 243238
rect 31760 242208 31812 242214
rect 31760 242150 31812 242156
rect 32404 241052 32456 241058
rect 32404 240994 32456 241000
rect 32416 189038 32444 240994
rect 32404 189032 32456 189038
rect 32404 188974 32456 188980
rect 32692 178022 32720 251874
rect 32772 242820 32824 242826
rect 32772 242762 32824 242768
rect 32680 178016 32732 178022
rect 32680 177958 32732 177964
rect 32784 125186 32812 242762
rect 32876 131102 32904 297366
rect 32956 242616 33008 242622
rect 32956 242558 33008 242564
rect 32864 131096 32916 131102
rect 32864 131038 32916 131044
rect 32772 125180 32824 125186
rect 32772 125122 32824 125128
rect 31668 69012 31720 69018
rect 31668 68954 31720 68960
rect 31576 60716 31628 60722
rect 31576 60658 31628 60664
rect 32968 46918 32996 242558
rect 32956 46912 33008 46918
rect 32956 46854 33008 46860
rect 21364 45552 21416 45558
rect 21364 45494 21416 45500
rect 33060 42770 33088 347822
rect 33796 246294 33824 500958
rect 34428 336048 34480 336054
rect 34428 335990 34480 335996
rect 34336 334620 34388 334626
rect 34336 334562 34388 334568
rect 34244 264240 34296 264246
rect 34244 264182 34296 264188
rect 33968 253224 34020 253230
rect 33968 253166 34020 253172
rect 33784 246288 33836 246294
rect 33784 246230 33836 246236
rect 33784 245064 33836 245070
rect 33784 245006 33836 245012
rect 33796 164218 33824 245006
rect 33980 169726 34008 253166
rect 34060 246628 34112 246634
rect 34060 246570 34112 246576
rect 33968 169720 34020 169726
rect 33968 169662 34020 169668
rect 33784 164212 33836 164218
rect 33784 164154 33836 164160
rect 34072 139398 34100 246570
rect 34152 241936 34204 241942
rect 34152 241878 34204 241884
rect 34060 139392 34112 139398
rect 34060 139334 34112 139340
rect 34164 121446 34192 241878
rect 34152 121440 34204 121446
rect 34152 121382 34204 121388
rect 34256 95198 34284 264182
rect 34348 161430 34376 334562
rect 34336 161424 34388 161430
rect 34336 161366 34388 161372
rect 34440 109002 34468 335990
rect 35072 246356 35124 246362
rect 35072 246298 35124 246304
rect 34428 108996 34480 109002
rect 34428 108938 34480 108944
rect 34244 95192 34296 95198
rect 34244 95134 34296 95140
rect 35084 56574 35112 246298
rect 35176 245342 35204 632062
rect 39672 425740 39724 425746
rect 39672 425682 39724 425688
rect 38474 376952 38530 376961
rect 38474 376887 38530 376896
rect 37922 376000 37978 376009
rect 37922 375935 37978 375944
rect 37830 348120 37886 348129
rect 37830 348055 37886 348064
rect 37844 347886 37872 348055
rect 37832 347880 37884 347886
rect 37832 347822 37884 347828
rect 35716 334688 35768 334694
rect 35716 334630 35768 334636
rect 35440 252136 35492 252142
rect 35440 252078 35492 252084
rect 35164 245336 35216 245342
rect 35164 245278 35216 245284
rect 35256 244928 35308 244934
rect 35256 244870 35308 244876
rect 35268 111790 35296 244870
rect 35348 242412 35400 242418
rect 35348 242354 35400 242360
rect 35360 195974 35388 242354
rect 35348 195968 35400 195974
rect 35348 195910 35400 195916
rect 35452 173398 35480 252078
rect 35532 242548 35584 242554
rect 35532 242490 35584 242496
rect 35440 173392 35492 173398
rect 35440 173334 35492 173340
rect 35544 151774 35572 242490
rect 35624 242004 35676 242010
rect 35624 241946 35676 241952
rect 35532 151768 35584 151774
rect 35532 151710 35584 151716
rect 35636 113150 35664 241946
rect 35728 147626 35756 334630
rect 37004 256012 37056 256018
rect 37004 255954 37056 255960
rect 35808 253632 35860 253638
rect 35808 253574 35860 253580
rect 35820 218006 35848 253574
rect 36912 250572 36964 250578
rect 36912 250514 36964 250520
rect 36728 249620 36780 249626
rect 36728 249562 36780 249568
rect 36636 243568 36688 243574
rect 36636 243510 36688 243516
rect 36544 242956 36596 242962
rect 36544 242898 36596 242904
rect 36452 242480 36504 242486
rect 36452 242422 36504 242428
rect 35808 218000 35860 218006
rect 35808 217942 35860 217948
rect 36464 187678 36492 242422
rect 36452 187672 36504 187678
rect 36452 187614 36504 187620
rect 35716 147620 35768 147626
rect 35716 147562 35768 147568
rect 35624 113144 35676 113150
rect 35624 113086 35676 113092
rect 35256 111784 35308 111790
rect 35256 111726 35308 111732
rect 35072 56568 35124 56574
rect 35072 56510 35124 56516
rect 33048 42764 33100 42770
rect 33048 42706 33100 42712
rect 36556 39370 36584 242898
rect 36648 213081 36676 243510
rect 36634 213072 36690 213081
rect 36634 213007 36690 213016
rect 36740 199889 36768 249562
rect 36820 246764 36872 246770
rect 36820 246706 36872 246712
rect 36726 199880 36782 199889
rect 36726 199815 36782 199824
rect 36832 164937 36860 246706
rect 36818 164928 36874 164937
rect 36818 164863 36874 164872
rect 36924 156097 36952 250514
rect 36910 156088 36966 156097
rect 36910 156023 36966 156032
rect 37016 143041 37044 255954
rect 37096 250980 37148 250986
rect 37096 250922 37148 250928
rect 37108 234977 37136 250922
rect 37188 242344 37240 242350
rect 37188 242286 37240 242292
rect 37094 234968 37150 234977
rect 37094 234903 37150 234912
rect 37200 226273 37228 242286
rect 37832 241392 37884 241398
rect 37832 241334 37884 241340
rect 37740 241120 37792 241126
rect 37740 241062 37792 241068
rect 37186 226264 37242 226273
rect 37186 226199 37242 226208
rect 37372 187672 37424 187678
rect 37372 187614 37424 187620
rect 37384 186833 37412 187614
rect 37370 186824 37426 186833
rect 37370 186759 37426 186768
rect 37096 186380 37148 186386
rect 37096 186322 37148 186328
rect 37002 143032 37058 143041
rect 37002 142967 37058 142976
rect 36544 39364 36596 39370
rect 36544 39306 36596 39312
rect 37108 38554 37136 186322
rect 37752 116657 37780 241062
rect 37844 221785 37872 241334
rect 37830 221776 37886 221785
rect 37830 221711 37886 221720
rect 37832 186448 37884 186454
rect 37832 186390 37884 186396
rect 37738 116648 37794 116657
rect 37738 116583 37794 116592
rect 37648 108996 37700 109002
rect 37648 108938 37700 108944
rect 37660 107953 37688 108938
rect 37646 107944 37702 107953
rect 37646 107879 37702 107888
rect 37844 50969 37872 186390
rect 37936 186386 37964 375935
rect 38106 373824 38162 373833
rect 38106 373759 38162 373768
rect 38120 339454 38148 373759
rect 38290 372872 38346 372881
rect 38290 372807 38346 372816
rect 38108 339448 38160 339454
rect 38108 339390 38160 339396
rect 38304 339386 38332 372807
rect 38382 350024 38438 350033
rect 38382 349959 38438 349968
rect 38292 339380 38344 339386
rect 38292 339322 38344 339328
rect 38108 247784 38160 247790
rect 38108 247726 38160 247732
rect 38016 218000 38068 218006
rect 38016 217942 38068 217948
rect 38028 217433 38056 217942
rect 38014 217424 38070 217433
rect 38014 217359 38070 217368
rect 38016 195968 38068 195974
rect 38016 195910 38068 195916
rect 38028 195537 38056 195910
rect 38014 195528 38070 195537
rect 38014 195463 38070 195472
rect 38016 191820 38068 191826
rect 38016 191762 38068 191768
rect 38028 191185 38056 191762
rect 38014 191176 38070 191185
rect 38014 191111 38070 191120
rect 37924 186380 37976 186386
rect 37924 186322 37976 186328
rect 38016 178016 38068 178022
rect 38014 177984 38016 177993
rect 38068 177984 38070 177993
rect 38014 177919 38070 177928
rect 38014 173632 38070 173641
rect 38014 173567 38070 173576
rect 38028 173398 38056 173567
rect 38016 173392 38068 173398
rect 38016 173334 38068 173340
rect 38016 169720 38068 169726
rect 38016 169662 38068 169668
rect 38028 169289 38056 169662
rect 38014 169280 38070 169289
rect 38014 169215 38070 169224
rect 38016 161424 38068 161430
rect 38016 161366 38068 161372
rect 38028 160449 38056 161366
rect 38014 160440 38070 160449
rect 38014 160375 38070 160384
rect 38016 151768 38068 151774
rect 38014 151736 38016 151745
rect 38068 151736 38070 151745
rect 38014 151671 38070 151680
rect 38016 147620 38068 147626
rect 38016 147562 38068 147568
rect 38028 147393 38056 147562
rect 38014 147384 38070 147393
rect 38014 147319 38070 147328
rect 38016 139392 38068 139398
rect 38016 139334 38068 139340
rect 38028 138553 38056 139334
rect 38014 138544 38070 138553
rect 38014 138479 38070 138488
rect 38120 134201 38148 247726
rect 38292 241324 38344 241330
rect 38292 241266 38344 241272
rect 38106 134192 38162 134201
rect 38106 134127 38162 134136
rect 38016 131096 38068 131102
rect 38016 131038 38068 131044
rect 38028 129849 38056 131038
rect 38014 129840 38070 129849
rect 38014 129775 38070 129784
rect 38014 125488 38070 125497
rect 38014 125423 38070 125432
rect 38028 125186 38056 125423
rect 38016 125180 38068 125186
rect 38016 125122 38068 125128
rect 37924 121440 37976 121446
rect 37924 121382 37976 121388
rect 37936 121009 37964 121382
rect 37922 121000 37978 121009
rect 37922 120935 37978 120944
rect 38200 117972 38252 117978
rect 38200 117914 38252 117920
rect 38016 113144 38068 113150
rect 38016 113086 38068 113092
rect 38028 112305 38056 113086
rect 38014 112296 38070 112305
rect 38014 112231 38070 112240
rect 38016 95192 38068 95198
rect 38016 95134 38068 95140
rect 38028 94761 38056 95134
rect 38014 94752 38070 94761
rect 38014 94687 38070 94696
rect 38016 91044 38068 91050
rect 38016 90986 38068 90992
rect 38028 90409 38056 90986
rect 38014 90400 38070 90409
rect 38014 90335 38070 90344
rect 38014 77208 38070 77217
rect 38014 77143 38070 77152
rect 38028 76974 38056 77143
rect 38016 76968 38068 76974
rect 38016 76910 38068 76916
rect 38016 69012 38068 69018
rect 38016 68954 38068 68960
rect 38028 68513 38056 68954
rect 38014 68504 38070 68513
rect 38014 68439 38070 68448
rect 38212 64161 38240 117914
rect 38304 99113 38332 241266
rect 38396 183530 38424 349959
rect 38384 183524 38436 183530
rect 38384 183466 38436 183472
rect 38290 99104 38346 99113
rect 38290 99039 38346 99048
rect 38198 64152 38254 64161
rect 38198 64087 38254 64096
rect 38016 60716 38068 60722
rect 38016 60658 38068 60664
rect 38028 59673 38056 60658
rect 38014 59664 38070 59673
rect 38014 59599 38070 59608
rect 38016 56568 38068 56574
rect 38016 56510 38068 56516
rect 38028 55321 38056 56510
rect 38014 55312 38070 55321
rect 38014 55247 38070 55256
rect 37830 50960 37886 50969
rect 37830 50895 37886 50904
rect 38016 46912 38068 46918
rect 38016 46854 38068 46860
rect 38028 46617 38056 46854
rect 38014 46608 38070 46617
rect 38014 46543 38070 46552
rect 38016 42764 38068 42770
rect 38016 42706 38068 42712
rect 38028 42265 38056 42706
rect 38014 42256 38070 42265
rect 38014 42191 38070 42200
rect 38488 38690 38516 376887
rect 38842 371104 38898 371113
rect 38842 371039 38898 371048
rect 38658 370016 38714 370025
rect 38658 369951 38714 369960
rect 38566 348392 38622 348401
rect 38566 348327 38622 348336
rect 38580 338094 38608 348327
rect 38568 338088 38620 338094
rect 38568 338030 38620 338036
rect 38580 242894 38608 338030
rect 38672 333402 38700 369951
rect 38750 368248 38806 368257
rect 38750 368183 38806 368192
rect 38660 333396 38712 333402
rect 38660 333338 38712 333344
rect 38660 324964 38712 324970
rect 38660 324906 38712 324912
rect 38568 242888 38620 242894
rect 38568 242830 38620 242836
rect 38568 241256 38620 241262
rect 38568 241198 38620 241204
rect 38580 86057 38608 241198
rect 38672 103601 38700 324906
rect 38764 278050 38792 368183
rect 38856 339046 38884 371039
rect 38844 339040 38896 339046
rect 38844 338982 38896 338988
rect 39396 337204 39448 337210
rect 39396 337146 39448 337152
rect 38752 278044 38804 278050
rect 38752 277986 38804 277992
rect 39304 242888 39356 242894
rect 39304 242830 39356 242836
rect 39212 242276 39264 242282
rect 39212 242218 39264 242224
rect 39028 242140 39080 242146
rect 39028 242082 39080 242088
rect 38844 241188 38896 241194
rect 38844 241130 38896 241136
rect 38752 240848 38804 240854
rect 38752 240790 38804 240796
rect 38658 103592 38714 103601
rect 38658 103527 38714 103536
rect 38566 86048 38622 86057
rect 38566 85983 38622 85992
rect 38764 72865 38792 240790
rect 38856 81569 38884 241130
rect 38936 240780 38988 240786
rect 38936 240722 38988 240728
rect 38948 182345 38976 240722
rect 39040 204377 39068 242082
rect 39120 241528 39172 241534
rect 39120 241470 39172 241476
rect 39132 208729 39160 241470
rect 39224 230625 39252 242218
rect 39210 230616 39266 230625
rect 39210 230551 39266 230560
rect 39118 208720 39174 208729
rect 39118 208655 39174 208664
rect 39026 204368 39082 204377
rect 39026 204303 39082 204312
rect 38934 182336 38990 182345
rect 38934 182271 38990 182280
rect 38842 81560 38898 81569
rect 38842 81495 38898 81504
rect 38750 72856 38806 72865
rect 38750 72791 38806 72800
rect 38476 38684 38528 38690
rect 38476 38626 38528 38632
rect 39316 38622 39344 242830
rect 39408 117978 39436 337146
rect 39684 243710 39712 425682
rect 39776 338706 39804 699654
rect 39764 338700 39816 338706
rect 39764 338642 39816 338648
rect 39672 243704 39724 243710
rect 39672 243646 39724 243652
rect 39868 243642 39896 700266
rect 40512 699718 40540 703520
rect 72988 699718 73016 703520
rect 89180 700330 89208 703520
rect 105464 700398 105492 703520
rect 105452 700392 105504 700398
rect 105452 700334 105504 700340
rect 106188 700392 106240 700398
rect 106188 700334 106240 700340
rect 89168 700324 89220 700330
rect 89168 700266 89220 700272
rect 40500 699712 40552 699718
rect 40500 699654 40552 699660
rect 71780 699712 71832 699718
rect 71780 699654 71832 699660
rect 72976 699712 73028 699718
rect 72976 699654 73028 699660
rect 71792 425746 71820 699654
rect 106200 425746 106228 700334
rect 137848 700330 137876 703520
rect 154132 702434 154160 703520
rect 153212 702406 154160 702434
rect 137836 700324 137888 700330
rect 137836 700266 137888 700272
rect 153212 474026 153240 702406
rect 170324 700398 170352 703520
rect 202800 703050 202828 703520
rect 201500 703044 201552 703050
rect 201500 702986 201552 702992
rect 202788 703044 202840 703050
rect 202788 702986 202840 702992
rect 170312 700392 170364 700398
rect 170312 700334 170364 700340
rect 178040 700392 178092 700398
rect 178040 700334 178092 700340
rect 193864 700392 193916 700398
rect 193864 700334 193916 700340
rect 176660 700324 176712 700330
rect 176660 700266 176712 700272
rect 153200 474020 153252 474026
rect 153200 473962 153252 473968
rect 71780 425740 71832 425746
rect 71780 425682 71832 425688
rect 106188 425740 106240 425746
rect 106188 425682 106240 425688
rect 131764 339448 131816 339454
rect 131764 339390 131816 339396
rect 92296 338972 92348 338978
rect 92296 338914 92348 338920
rect 81348 338904 81400 338910
rect 81348 338846 81400 338852
rect 75828 338836 75880 338842
rect 75828 338778 75880 338784
rect 73068 338768 73120 338774
rect 73068 338710 73120 338716
rect 48964 338020 49016 338026
rect 48964 337962 49016 337968
rect 40500 337952 40552 337958
rect 40500 337894 40552 337900
rect 40408 337272 40460 337278
rect 40408 337214 40460 337220
rect 39856 243636 39908 243642
rect 39856 243578 39908 243584
rect 39856 242888 39908 242894
rect 39856 242830 39908 242836
rect 39868 241534 39896 242830
rect 39948 242072 40000 242078
rect 39948 242014 40000 242020
rect 39856 241528 39908 241534
rect 39856 241470 39908 241476
rect 39960 239873 39988 242014
rect 39946 239864 40002 239873
rect 39946 239799 40002 239808
rect 39488 183524 39540 183530
rect 39488 183466 39540 183472
rect 39396 117972 39448 117978
rect 39396 117914 39448 117920
rect 39304 38616 39356 38622
rect 39304 38558 39356 38564
rect 37096 38548 37148 38554
rect 37096 38490 37148 38496
rect 39500 38418 39528 183466
rect 40420 38486 40448 337214
rect 40512 186454 40540 337894
rect 43444 337816 43496 337822
rect 43444 337758 43496 337764
rect 42064 337000 42116 337006
rect 42064 336942 42116 336948
rect 41786 244352 41842 244361
rect 41786 244287 41842 244296
rect 40592 242956 40644 242962
rect 40592 242898 40644 242904
rect 40604 241468 40632 242898
rect 41800 241468 41828 244287
rect 42076 241262 42104 336942
rect 43456 241398 43484 337758
rect 48044 244452 48096 244458
rect 48044 244394 48096 244400
rect 44272 244384 44324 244390
rect 44272 244326 44324 244332
rect 44284 241468 44312 244326
rect 46848 243364 46900 243370
rect 46848 243306 46900 243312
rect 46860 241468 46888 243306
rect 48056 241468 48084 244394
rect 43444 241392 43496 241398
rect 43444 241334 43496 241340
rect 48976 241330 49004 337962
rect 56506 337920 56562 337929
rect 56506 337855 56508 337864
rect 56560 337855 56562 337864
rect 56508 337826 56560 337832
rect 68926 337784 68982 337793
rect 68926 337719 68982 337728
rect 70582 337784 70638 337793
rect 70582 337719 70638 337728
rect 59266 337648 59322 337657
rect 59266 337583 59322 337592
rect 62026 337648 62082 337657
rect 62026 337583 62082 337592
rect 63406 337648 63462 337657
rect 63406 337583 63462 337592
rect 64970 337648 65026 337657
rect 64970 337583 65026 337592
rect 66350 337648 66406 337657
rect 66350 337583 66406 337592
rect 67638 337648 67694 337657
rect 67638 337583 67694 337592
rect 57886 337512 57942 337521
rect 57886 337447 57942 337456
rect 57900 337414 57928 337447
rect 57888 337408 57940 337414
rect 57888 337350 57940 337356
rect 50344 336864 50396 336870
rect 50344 336806 50396 336812
rect 48964 241324 49016 241330
rect 48964 241266 49016 241272
rect 50356 241262 50384 336806
rect 59280 247926 59308 337583
rect 59450 337376 59506 337385
rect 59450 337311 59506 337320
rect 59464 337278 59492 337311
rect 59452 337272 59504 337278
rect 59358 337240 59414 337249
rect 59452 337214 59504 337220
rect 59358 337175 59360 337184
rect 59412 337175 59414 337184
rect 59360 337146 59412 337152
rect 59268 247920 59320 247926
rect 59268 247862 59320 247868
rect 62040 247858 62068 337583
rect 62028 247852 62080 247858
rect 62028 247794 62080 247800
rect 59360 244656 59412 244662
rect 59360 244598 59412 244604
rect 55588 244588 55640 244594
rect 55588 244530 55640 244536
rect 51816 244520 51868 244526
rect 51816 244462 51868 244468
rect 51828 241468 51856 244462
rect 55600 241468 55628 244530
rect 58072 243228 58124 243234
rect 58072 243170 58124 243176
rect 58084 241468 58112 243170
rect 59372 241468 59400 244598
rect 63132 243772 63184 243778
rect 63132 243714 63184 243720
rect 60648 243500 60700 243506
rect 60648 243442 60700 243448
rect 60660 241468 60688 243442
rect 61844 243432 61896 243438
rect 61844 243374 61896 243380
rect 61856 241468 61884 243374
rect 63144 241468 63172 243714
rect 63420 242690 63448 337583
rect 64786 337512 64842 337521
rect 64786 337447 64842 337456
rect 64696 271924 64748 271930
rect 64696 271866 64748 271872
rect 63408 242684 63460 242690
rect 63408 242626 63460 242632
rect 64708 241482 64736 271866
rect 64800 242214 64828 337447
rect 64788 242208 64840 242214
rect 64788 242150 64840 242156
rect 64446 241454 64736 241482
rect 42064 241256 42116 241262
rect 50344 241256 50396 241262
rect 42064 241198 42116 241204
rect 45586 241194 45968 241210
rect 49358 241194 49648 241210
rect 57152 241256 57204 241262
rect 50344 241198 50396 241204
rect 50646 241194 50936 241210
rect 53130 241194 53512 241210
rect 54326 241194 54616 241210
rect 56902 241204 57152 241210
rect 56902 241198 57204 241204
rect 45586 241188 45980 241194
rect 45586 241182 45928 241188
rect 49358 241188 49660 241194
rect 49358 241182 49608 241188
rect 45928 241130 45980 241136
rect 50646 241188 50948 241194
rect 50646 241182 50896 241188
rect 49608 241130 49660 241136
rect 53130 241188 53524 241194
rect 53130 241182 53472 241188
rect 50896 241130 50948 241136
rect 54326 241188 54628 241194
rect 54326 241182 54576 241188
rect 53472 241130 53524 241136
rect 56902 241182 57192 241198
rect 64984 241194 65012 337583
rect 66168 258120 66220 258126
rect 66168 258062 66220 258068
rect 66180 248414 66208 258062
rect 66088 248386 66208 248414
rect 66088 241482 66116 248386
rect 65642 241454 66116 241482
rect 64972 241188 65024 241194
rect 54576 241130 54628 241136
rect 64972 241130 65024 241136
rect 66364 241126 66392 337583
rect 67652 324970 67680 337583
rect 67640 324964 67692 324970
rect 67640 324906 67692 324912
rect 68836 324352 68888 324358
rect 68836 324294 68888 324300
rect 67548 298172 67600 298178
rect 67548 298114 67600 298120
rect 67560 248414 67588 298114
rect 67376 248386 67588 248414
rect 67376 241482 67404 248386
rect 68848 244254 68876 324294
rect 68100 244248 68152 244254
rect 68100 244190 68152 244196
rect 68836 244248 68888 244254
rect 68836 244190 68888 244196
rect 66930 241454 67404 241482
rect 68112 241468 68140 244190
rect 68940 242758 68968 337719
rect 70490 337648 70546 337657
rect 70490 337583 70546 337592
rect 69110 337376 69166 337385
rect 69110 337311 69166 337320
rect 68928 242752 68980 242758
rect 68928 242694 68980 242700
rect 69124 241942 69152 337311
rect 70308 311908 70360 311914
rect 70308 311850 70360 311856
rect 70320 244254 70348 311850
rect 70504 246362 70532 337583
rect 70492 246356 70544 246362
rect 70492 246298 70544 246304
rect 69388 244248 69440 244254
rect 69388 244190 69440 244196
rect 70308 244248 70360 244254
rect 70308 244190 70360 244196
rect 69112 241936 69164 241942
rect 69112 241878 69164 241884
rect 69400 241468 69428 244190
rect 70596 242826 70624 337719
rect 72974 337512 73030 337521
rect 72974 337447 73030 337456
rect 72988 337278 73016 337447
rect 72976 337272 73028 337278
rect 72976 337214 73028 337220
rect 71688 257372 71740 257378
rect 71688 257314 71740 257320
rect 71700 244254 71728 257314
rect 73080 244254 73108 338710
rect 74354 337784 74410 337793
rect 74354 337719 74410 337728
rect 74368 254590 74396 337719
rect 74446 337648 74502 337657
rect 74446 337583 74502 337592
rect 74906 337648 74962 337657
rect 74906 337583 74962 337592
rect 74356 254584 74408 254590
rect 74356 254526 74408 254532
rect 74460 252074 74488 337583
rect 74920 334898 74948 337583
rect 74908 334892 74960 334898
rect 74908 334834 74960 334840
rect 74448 252068 74500 252074
rect 74448 252010 74500 252016
rect 74448 250504 74500 250510
rect 74448 250446 74500 250452
rect 73160 246424 73212 246430
rect 73160 246366 73212 246372
rect 70676 244248 70728 244254
rect 70676 244190 70728 244196
rect 71688 244248 71740 244254
rect 71688 244190 71740 244196
rect 71872 244248 71924 244254
rect 71872 244190 71924 244196
rect 73068 244248 73120 244254
rect 73068 244190 73120 244196
rect 70584 242820 70636 242826
rect 70584 242762 70636 242768
rect 70688 241468 70716 244190
rect 71884 241468 71912 244190
rect 73172 241468 73200 246366
rect 74460 241468 74488 250446
rect 75840 241482 75868 338778
rect 76286 338056 76342 338065
rect 76286 337991 76342 338000
rect 76300 334830 76328 337991
rect 78586 337920 78642 337929
rect 78586 337855 78642 337864
rect 77206 337784 77262 337793
rect 77206 337719 77262 337728
rect 77220 337482 77248 337719
rect 78494 337648 78550 337657
rect 78494 337583 78550 337592
rect 77208 337476 77260 337482
rect 77208 337418 77260 337424
rect 77206 336832 77262 336841
rect 77206 336767 77262 336776
rect 77220 336190 77248 336767
rect 77208 336184 77260 336190
rect 77208 336126 77260 336132
rect 76288 334824 76340 334830
rect 76288 334766 76340 334772
rect 78508 254658 78536 337583
rect 78600 337550 78628 337855
rect 79966 337648 80022 337657
rect 79966 337583 80022 337592
rect 81070 337648 81126 337657
rect 81070 337583 81126 337592
rect 78588 337544 78640 337550
rect 78588 337486 78640 337492
rect 79980 269822 80008 337583
rect 81084 334966 81112 337583
rect 81254 336832 81310 336841
rect 81254 336767 81310 336776
rect 81268 336326 81296 336767
rect 81256 336320 81308 336326
rect 81256 336262 81308 336268
rect 81072 334960 81124 334966
rect 81072 334902 81124 334908
rect 79968 269816 80020 269822
rect 79968 269758 80020 269764
rect 78496 254652 78548 254658
rect 78496 254594 78548 254600
rect 79416 250912 79468 250918
rect 79416 250854 79468 250860
rect 78220 249484 78272 249490
rect 78220 249426 78272 249432
rect 76932 246492 76984 246498
rect 76932 246434 76984 246440
rect 75670 241454 75868 241482
rect 76944 241468 76972 246434
rect 78232 241468 78260 249426
rect 79428 241468 79456 250854
rect 81360 248414 81388 338846
rect 91006 338056 91062 338065
rect 91006 337991 91062 338000
rect 83554 337784 83610 337793
rect 83554 337719 83610 337728
rect 88062 337784 88118 337793
rect 88062 337719 88118 337728
rect 82726 337648 82782 337657
rect 82726 337583 82782 337592
rect 82910 337648 82966 337657
rect 82910 337583 82966 337592
rect 81900 250640 81952 250646
rect 81900 250582 81952 250588
rect 81176 248386 81388 248414
rect 81176 241482 81204 248386
rect 80730 241454 81204 241482
rect 81912 241468 81940 250582
rect 82740 242826 82768 337583
rect 82728 242820 82780 242826
rect 82728 242762 82780 242768
rect 82924 242010 82952 337583
rect 83002 336968 83058 336977
rect 83002 336903 83058 336912
rect 82912 242004 82964 242010
rect 82912 241946 82964 241952
rect 83016 241126 83044 336903
rect 83568 333334 83596 337719
rect 85302 337648 85358 337657
rect 85302 337583 85358 337592
rect 86406 337648 86462 337657
rect 86406 337583 86462 337592
rect 85316 333606 85344 337583
rect 85304 333600 85356 333606
rect 85304 333542 85356 333548
rect 86420 333538 86448 337583
rect 86408 333532 86460 333538
rect 86408 333474 86460 333480
rect 83556 333328 83608 333334
rect 83556 333270 83608 333276
rect 85488 262880 85540 262886
rect 85488 262822 85540 262828
rect 83188 249416 83240 249422
rect 83188 249358 83240 249364
rect 83200 241468 83228 249358
rect 85500 244254 85528 262822
rect 85672 249076 85724 249082
rect 85672 249018 85724 249024
rect 84476 244248 84528 244254
rect 84476 244190 84528 244196
rect 85488 244248 85540 244254
rect 85488 244190 85540 244196
rect 84488 241468 84516 244190
rect 85684 241468 85712 249018
rect 86960 244248 87012 244254
rect 86960 244190 87012 244196
rect 86972 241468 87000 244190
rect 88076 241126 88104 337719
rect 88154 337648 88210 337657
rect 88154 337583 88210 337592
rect 88430 337648 88486 337657
rect 88430 337583 88486 337592
rect 90638 337648 90694 337657
rect 91020 337618 91048 337991
rect 91190 337648 91246 337657
rect 90638 337583 90694 337592
rect 91008 337612 91060 337618
rect 88168 268394 88196 337583
rect 88156 268388 88208 268394
rect 88156 268330 88208 268336
rect 88156 260160 88208 260166
rect 88156 260102 88208 260108
rect 88168 244254 88196 260102
rect 88248 246968 88300 246974
rect 88248 246910 88300 246916
rect 88156 244248 88208 244254
rect 88156 244190 88208 244196
rect 88260 241468 88288 246910
rect 88444 242146 88472 337583
rect 90652 333470 90680 337583
rect 91190 337583 91246 337592
rect 91008 337554 91060 337560
rect 90640 333464 90692 333470
rect 90640 333406 90692 333412
rect 90732 251048 90784 251054
rect 90732 250990 90784 250996
rect 89444 249688 89496 249694
rect 89444 249630 89496 249636
rect 88432 242140 88484 242146
rect 88432 242082 88484 242088
rect 89456 241468 89484 249630
rect 90744 241468 90772 250990
rect 91204 242894 91232 337583
rect 91192 242888 91244 242894
rect 91192 242830 91244 242836
rect 92308 241482 92336 338914
rect 126980 338700 127032 338706
rect 126980 338642 127032 338648
rect 99286 337920 99342 337929
rect 99286 337855 99342 337864
rect 92386 337784 92442 337793
rect 92386 337719 92442 337728
rect 93582 337784 93638 337793
rect 93582 337719 93638 337728
rect 95146 337784 95202 337793
rect 95146 337719 95202 337728
rect 97998 337784 98054 337793
rect 99300 337754 99328 337855
rect 97998 337719 98054 337728
rect 99288 337748 99340 337754
rect 92400 242894 92428 337719
rect 92478 337648 92534 337657
rect 92478 337583 92534 337592
rect 92492 256018 92520 337583
rect 93596 336802 93624 337719
rect 95160 337686 95188 337719
rect 95148 337680 95200 337686
rect 95148 337622 95200 337628
rect 96342 337648 96398 337657
rect 96342 337583 96398 337592
rect 97906 337648 97962 337657
rect 97906 337583 97962 337592
rect 93584 336796 93636 336802
rect 93584 336738 93636 336744
rect 92480 256012 92532 256018
rect 92480 255954 92532 255960
rect 93216 249756 93268 249762
rect 93216 249698 93268 249704
rect 92388 242888 92440 242894
rect 92388 242830 92440 242836
rect 92046 241454 92336 241482
rect 93228 241468 93256 249698
rect 94504 249552 94556 249558
rect 94504 249494 94556 249500
rect 94516 241468 94544 249494
rect 95700 247036 95752 247042
rect 95700 246978 95752 246984
rect 95712 241468 95740 246978
rect 96356 242146 96384 337583
rect 96526 336832 96582 336841
rect 96526 336767 96582 336776
rect 96540 336462 96568 336767
rect 96528 336456 96580 336462
rect 96528 336398 96580 336404
rect 97920 273970 97948 337583
rect 97908 273964 97960 273970
rect 97908 273906 97960 273912
rect 96988 249144 97040 249150
rect 96988 249086 97040 249092
rect 96344 242140 96396 242146
rect 96344 242082 96396 242088
rect 97000 241468 97028 249086
rect 98012 242078 98040 337719
rect 99288 337690 99340 337696
rect 100758 337648 100814 337657
rect 100758 337583 100814 337592
rect 106186 337648 106242 337657
rect 106186 337583 106242 337592
rect 107658 337648 107714 337657
rect 107658 337583 107714 337592
rect 111706 337648 111762 337657
rect 111706 337583 111762 337592
rect 113178 337648 113234 337657
rect 113178 337583 113234 337592
rect 118606 337648 118662 337657
rect 118606 337583 118662 337592
rect 121366 337648 121422 337657
rect 121366 337583 121422 337592
rect 122838 337648 122894 337657
rect 122838 337583 122894 337592
rect 126886 337648 126942 337657
rect 126886 337583 126942 337592
rect 99286 336832 99342 336841
rect 99286 336767 99342 336776
rect 100024 336796 100076 336802
rect 99300 336530 99328 336767
rect 100024 336738 100076 336744
rect 99288 336524 99340 336530
rect 99288 336466 99340 336472
rect 100036 271182 100064 336738
rect 100024 271176 100076 271182
rect 100024 271118 100076 271124
rect 100024 261520 100076 261526
rect 100024 261462 100076 261468
rect 99472 246356 99524 246362
rect 99472 246298 99524 246304
rect 98276 244248 98328 244254
rect 98276 244190 98328 244196
rect 98000 242072 98052 242078
rect 98000 242014 98052 242020
rect 98288 241468 98316 244190
rect 99484 241468 99512 246298
rect 100036 244254 100064 261462
rect 100772 250578 100800 337583
rect 104806 336832 104862 336841
rect 104806 336767 104862 336776
rect 104716 253360 104768 253366
rect 104716 253302 104768 253308
rect 102048 251864 102100 251870
rect 102048 251806 102100 251812
rect 100760 250572 100812 250578
rect 100760 250514 100812 250520
rect 101956 250572 102008 250578
rect 101956 250514 102008 250520
rect 100760 244316 100812 244322
rect 100760 244258 100812 244264
rect 100024 244248 100076 244254
rect 100024 244190 100076 244196
rect 100772 243778 100800 244258
rect 100760 243772 100812 243778
rect 100760 243714 100812 243720
rect 100760 242956 100812 242962
rect 100760 242898 100812 242904
rect 100772 241468 100800 242898
rect 101968 241482 101996 250514
rect 102060 242962 102088 251806
rect 103244 246560 103296 246566
rect 103244 246502 103296 246508
rect 102048 242956 102100 242962
rect 102048 242898 102100 242904
rect 101968 241454 102074 241482
rect 103256 241468 103284 246502
rect 104728 241482 104756 253302
rect 104820 249286 104848 336767
rect 106096 252000 106148 252006
rect 106096 251942 106148 251948
rect 104808 249280 104860 249286
rect 104808 249222 104860 249228
rect 106108 241482 106136 251942
rect 106200 250714 106228 337583
rect 107568 264308 107620 264314
rect 107568 264250 107620 264256
rect 106188 250708 106240 250714
rect 106188 250650 106240 250656
rect 107580 248414 107608 264250
rect 107488 248386 107608 248414
rect 107488 241482 107516 248386
rect 107672 246770 107700 337583
rect 108764 256012 108816 256018
rect 108764 255954 108816 255960
rect 107660 246764 107712 246770
rect 107660 246706 107712 246712
rect 108776 241482 108804 255954
rect 111616 252340 111668 252346
rect 111616 252282 111668 252288
rect 109500 251116 109552 251122
rect 109500 251058 109552 251064
rect 104558 241454 104756 241482
rect 105846 241454 106136 241482
rect 107042 241454 107516 241482
rect 108330 241454 108804 241482
rect 109512 241468 109540 251058
rect 111628 244254 111656 252282
rect 111720 246838 111748 337583
rect 113192 252142 113220 337583
rect 117226 337240 117282 337249
rect 117226 337175 117282 337184
rect 117240 336258 117268 337175
rect 117228 336252 117280 336258
rect 117228 336194 117280 336200
rect 118620 253570 118648 337583
rect 119988 336592 120040 336598
rect 119988 336534 120040 336540
rect 118608 253564 118660 253570
rect 118608 253506 118660 253512
rect 117964 252408 118016 252414
rect 117964 252350 118016 252356
rect 113180 252136 113232 252142
rect 113180 252078 113232 252084
rect 114468 252136 114520 252142
rect 114468 252078 114520 252084
rect 111708 246832 111760 246838
rect 111708 246774 111760 246780
rect 112076 244996 112128 245002
rect 112076 244938 112128 244944
rect 110788 244248 110840 244254
rect 110788 244190 110840 244196
rect 111616 244248 111668 244254
rect 111616 244190 111668 244196
rect 110800 241468 110828 244190
rect 112088 241468 112116 244938
rect 114480 244254 114508 252078
rect 114560 246764 114612 246770
rect 114560 246706 114612 246712
rect 113272 244248 113324 244254
rect 113272 244190 113324 244196
rect 114468 244248 114520 244254
rect 114468 244190 114520 244196
rect 113284 241468 113312 244190
rect 114572 241468 114600 246706
rect 115848 245200 115900 245206
rect 115848 245142 115900 245148
rect 115860 241468 115888 245142
rect 117976 244254 118004 252350
rect 118332 246152 118384 246158
rect 118332 246094 118384 246100
rect 117044 244248 117096 244254
rect 117044 244190 117096 244196
rect 117964 244248 118016 244254
rect 117964 244190 118016 244196
rect 115940 243500 115992 243506
rect 115940 243442 115992 243448
rect 115952 241194 115980 243442
rect 117056 241468 117084 244190
rect 118344 241468 118372 246094
rect 120000 241482 120028 336534
rect 121380 249354 121408 337583
rect 122852 249626 122880 337583
rect 126900 265674 126928 337583
rect 126888 265668 126940 265674
rect 126888 265610 126940 265616
rect 122840 249620 122892 249626
rect 122840 249562 122892 249568
rect 121368 249348 121420 249354
rect 121368 249290 121420 249296
rect 123300 243908 123352 243914
rect 123300 243850 123352 243856
rect 122104 243840 122156 243846
rect 122104 243782 122156 243788
rect 120816 243772 120868 243778
rect 120816 243714 120868 243720
rect 119646 241454 120028 241482
rect 120828 241468 120856 243714
rect 122116 241468 122144 243782
rect 123312 241468 123340 243850
rect 124588 243704 124640 243710
rect 124588 243646 124640 243652
rect 124600 241468 124628 243646
rect 125876 243636 125928 243642
rect 125876 243578 125928 243584
rect 125888 241468 125916 243578
rect 126992 241482 127020 338642
rect 131026 338056 131082 338065
rect 131026 337991 131082 338000
rect 129646 337648 129702 337657
rect 129646 337583 129702 337592
rect 129660 253502 129688 337583
rect 131040 336394 131068 337991
rect 131028 336388 131080 336394
rect 131028 336330 131080 336336
rect 129648 253496 129700 253502
rect 129648 253438 129700 253444
rect 130844 249212 130896 249218
rect 130844 249154 130896 249160
rect 128360 246900 128412 246906
rect 128360 246842 128412 246848
rect 126992 241454 127098 241482
rect 128372 241468 128400 246842
rect 129648 246220 129700 246226
rect 129648 246162 129700 246168
rect 129660 241468 129688 246162
rect 130856 241468 130884 249154
rect 131776 243710 131804 339390
rect 153844 339380 153896 339386
rect 153844 339322 153896 339328
rect 132500 339312 132552 339318
rect 132500 339254 132552 339260
rect 132132 250844 132184 250850
rect 132132 250786 132184 250792
rect 131764 243704 131816 243710
rect 131764 243646 131816 243652
rect 132144 241468 132172 250786
rect 132512 241548 132540 339254
rect 136640 339244 136692 339250
rect 136640 339186 136692 339192
rect 132590 337648 132646 337657
rect 132590 337583 132646 337592
rect 135258 337648 135314 337657
rect 135258 337583 135314 337592
rect 132604 243574 132632 337583
rect 135272 253638 135300 337583
rect 135260 253632 135312 253638
rect 135260 253574 135312 253580
rect 135536 252272 135588 252278
rect 135536 252214 135588 252220
rect 134616 245336 134668 245342
rect 134616 245278 134668 245284
rect 132592 243568 132644 243574
rect 132592 243510 132644 243516
rect 132512 241520 133000 241548
rect 132972 241482 133000 241520
rect 132972 241454 133446 241482
rect 134628 241468 134656 245278
rect 135548 241482 135576 252214
rect 136652 241482 136680 339186
rect 140780 339176 140832 339182
rect 140780 339118 140832 339124
rect 139306 337648 139362 337657
rect 139306 337583 139362 337592
rect 139320 246906 139348 337583
rect 139400 282192 139452 282198
rect 139400 282134 139452 282140
rect 139308 246900 139360 246906
rect 139308 246842 139360 246848
rect 138388 245268 138440 245274
rect 138388 245210 138440 245216
rect 135548 241454 135930 241482
rect 136652 241454 137126 241482
rect 138400 241468 138428 245210
rect 139412 241482 139440 282134
rect 140792 241482 140820 339118
rect 142158 337784 142214 337793
rect 142158 337719 142214 337728
rect 142066 337648 142122 337657
rect 142066 337583 142122 337592
rect 142080 250850 142108 337583
rect 142172 250986 142200 337719
rect 146206 337648 146262 337657
rect 146206 337583 146262 337592
rect 143540 336116 143592 336122
rect 143540 336058 143592 336064
rect 143552 267734 143580 336058
rect 143552 267706 144224 267734
rect 142160 250980 142212 250986
rect 142160 250922 142212 250928
rect 142068 250844 142120 250850
rect 142068 250786 142120 250792
rect 142160 250776 142212 250782
rect 142160 250718 142212 250724
rect 139412 241454 139702 241482
rect 140792 241454 140898 241482
rect 142172 241468 142200 250718
rect 143448 246288 143500 246294
rect 143448 246230 143500 246236
rect 143460 241468 143488 246230
rect 144196 241482 144224 267706
rect 146220 249626 146248 337583
rect 150440 311160 150492 311166
rect 150440 311102 150492 311108
rect 146300 290488 146352 290494
rect 146300 290430 146352 290436
rect 146312 267734 146340 290430
rect 149060 280832 149112 280838
rect 149060 280774 149112 280780
rect 149072 267734 149100 280774
rect 146312 267706 146800 267734
rect 149072 267706 149376 267734
rect 146208 249620 146260 249626
rect 146208 249562 146260 249568
rect 145932 245132 145984 245138
rect 145932 245074 145984 245080
rect 144196 241454 144670 241482
rect 145944 241468 145972 245074
rect 146772 241482 146800 267706
rect 148048 253428 148100 253434
rect 148048 253370 148100 253376
rect 148060 241482 148088 253370
rect 149348 241482 149376 267706
rect 150452 241482 150480 311102
rect 153200 252204 153252 252210
rect 153200 252146 153252 252152
rect 152188 246696 152240 246702
rect 152188 246638 152240 246644
rect 146772 241454 147154 241482
rect 148060 241454 148442 241482
rect 149348 241454 149730 241482
rect 150452 241454 150926 241482
rect 152200 241468 152228 246638
rect 153212 241482 153240 252146
rect 153856 243982 153884 339322
rect 155960 339108 156012 339114
rect 155960 339050 156012 339056
rect 154580 260228 154632 260234
rect 154580 260170 154632 260176
rect 153844 243976 153896 243982
rect 153844 243918 153896 243924
rect 154592 241482 154620 260170
rect 153212 241454 153502 241482
rect 154592 241454 154698 241482
rect 155972 241468 156000 339050
rect 171784 336524 171836 336530
rect 171784 336466 171836 336472
rect 162124 333600 162176 333606
rect 162124 333542 162176 333548
rect 156052 318844 156104 318850
rect 156052 318786 156104 318792
rect 156064 267734 156092 318786
rect 158720 305040 158772 305046
rect 158720 304982 158772 304988
rect 157340 292596 157392 292602
rect 157340 292538 157392 292544
rect 157352 267734 157380 292538
rect 158732 267734 158760 304982
rect 156064 267706 156920 267734
rect 157352 267706 158024 267734
rect 158732 267706 159312 267734
rect 156892 241482 156920 267706
rect 157996 241482 158024 267706
rect 159284 241482 159312 267706
rect 160560 266416 160612 266422
rect 160560 266358 160612 266364
rect 160572 241482 160600 266358
rect 162136 244050 162164 333542
rect 169024 333532 169076 333538
rect 169024 333474 169076 333480
rect 167644 268388 167696 268394
rect 167644 268330 167696 268336
rect 163136 253972 163188 253978
rect 163136 253914 163188 253920
rect 162124 244044 162176 244050
rect 162124 243986 162176 243992
rect 162216 243296 162268 243302
rect 162216 243238 162268 243244
rect 156892 241454 157274 241482
rect 157996 241454 158470 241482
rect 159284 241454 159758 241482
rect 160572 241454 160954 241482
rect 162228 241468 162256 243238
rect 163148 241482 163176 253914
rect 164700 244860 164752 244866
rect 164700 244802 164752 244808
rect 163148 241454 163530 241482
rect 164712 241468 164740 244802
rect 167656 243506 167684 268330
rect 168472 245064 168524 245070
rect 168472 245006 168524 245012
rect 167644 243500 167696 243506
rect 167644 243442 167696 243448
rect 167276 243160 167328 243166
rect 167276 243102 167328 243108
rect 167288 241468 167316 243102
rect 168484 241468 168512 245006
rect 169036 244118 169064 333474
rect 171796 244186 171824 336466
rect 173164 336456 173216 336462
rect 173164 336398 173216 336404
rect 172244 244928 172296 244934
rect 172244 244870 172296 244876
rect 171048 244180 171100 244186
rect 171048 244122 171100 244128
rect 171784 244180 171836 244186
rect 171784 244122 171836 244128
rect 169024 244112 169076 244118
rect 169024 244054 169076 244060
rect 171060 241468 171088 244122
rect 172256 241468 172284 244870
rect 173176 244254 173204 336398
rect 176016 244792 176068 244798
rect 176016 244734 176068 244740
rect 173164 244248 173216 244254
rect 173164 244190 173216 244196
rect 172428 243364 172480 243370
rect 172428 243306 172480 243312
rect 115940 241188 115992 241194
rect 115940 241130 115992 241136
rect 43352 241120 43404 241126
rect 43102 241068 43352 241074
rect 43102 241062 43404 241068
rect 66352 241120 66404 241126
rect 66352 241062 66404 241068
rect 83004 241120 83056 241126
rect 83004 241062 83056 241068
rect 88064 241120 88116 241126
rect 88064 241062 88116 241068
rect 43102 241046 43392 241062
rect 165632 241058 166014 241074
rect 165620 241052 166014 241058
rect 165672 241046 166014 241052
rect 165620 240994 165672 241000
rect 172440 240990 172468 243306
rect 174728 243092 174780 243098
rect 174728 243034 174780 243040
rect 173176 241466 173558 241482
rect 174740 241468 174768 243034
rect 176028 241468 176056 244734
rect 176672 243778 176700 700266
rect 176752 474020 176804 474026
rect 176752 473962 176804 473968
rect 176764 243846 176792 473962
rect 176844 425740 176896 425746
rect 176844 425682 176896 425688
rect 176856 243914 176884 425682
rect 178052 336598 178080 700334
rect 191104 696992 191156 696998
rect 191104 696934 191156 696940
rect 182824 670744 182876 670750
rect 182824 670686 182876 670692
rect 180064 616888 180116 616894
rect 180064 616830 180116 616836
rect 178684 456816 178736 456822
rect 178684 456758 178736 456764
rect 178040 336592 178092 336598
rect 178040 336534 178092 336540
rect 177304 336320 177356 336326
rect 177304 336262 177356 336268
rect 176844 243908 176896 243914
rect 176844 243850 176896 243856
rect 176752 243840 176804 243846
rect 176752 243782 176804 243788
rect 177316 243778 177344 336262
rect 178696 249490 178724 456758
rect 180076 249694 180104 616830
rect 182836 249762 182864 670686
rect 189724 643136 189776 643142
rect 189724 643078 189776 643084
rect 186964 536852 187016 536858
rect 186964 536794 187016 536800
rect 185584 484424 185636 484430
rect 185584 484366 185636 484372
rect 184848 349172 184900 349178
rect 184848 349114 184900 349120
rect 182824 249756 182876 249762
rect 182824 249698 182876 249704
rect 180064 249688 180116 249694
rect 180064 249630 180116 249636
rect 178684 249484 178736 249490
rect 178684 249426 178736 249432
rect 179788 244724 179840 244730
rect 179788 244666 179840 244672
rect 176660 243772 176712 243778
rect 176660 243714 176712 243720
rect 177304 243772 177356 243778
rect 177304 243714 177356 243720
rect 178500 243024 178552 243030
rect 178500 242966 178552 242972
rect 178512 241468 178540 242966
rect 179800 241468 179828 244666
rect 184664 243432 184716 243438
rect 184664 243374 184716 243380
rect 183560 243364 183612 243370
rect 183560 243306 183612 243312
rect 183572 241468 183600 243306
rect 173164 241460 173558 241466
rect 173216 241454 173558 241460
rect 173164 241402 173216 241408
rect 169576 240984 169628 240990
rect 172428 240984 172480 240990
rect 169628 240932 169786 240938
rect 169576 240926 169786 240932
rect 172428 240926 172480 240932
rect 169588 240910 169786 240926
rect 177040 240922 177330 240938
rect 180904 240922 181102 240938
rect 182100 240922 182298 240938
rect 184676 240922 184704 243374
rect 184860 243370 184888 349114
rect 185596 250918 185624 484366
rect 185584 250912 185636 250918
rect 185584 250854 185636 250860
rect 186976 249422 187004 536794
rect 189080 333396 189132 333402
rect 189080 333338 189132 333344
rect 189092 267734 189120 333338
rect 189092 267706 189488 267734
rect 186964 249416 187016 249422
rect 186964 249358 187016 249364
rect 187332 247920 187384 247926
rect 187332 247862 187384 247868
rect 186044 243568 186096 243574
rect 186044 243510 186096 243516
rect 184848 243364 184900 243370
rect 184848 243306 184900 243312
rect 184846 242992 184902 243001
rect 184846 242927 184902 242936
rect 184860 241468 184888 242927
rect 186056 241468 186084 243510
rect 187344 241468 187372 247862
rect 188528 243636 188580 243642
rect 188528 243578 188580 243584
rect 187700 243228 187752 243234
rect 187700 243170 187752 243176
rect 187712 240990 187740 243170
rect 188540 241468 188568 243578
rect 189460 241482 189488 267706
rect 189736 251054 189764 643078
rect 189724 251048 189776 251054
rect 189724 250990 189776 250996
rect 191116 249558 191144 696934
rect 193128 369912 193180 369918
rect 193128 369854 193180 369860
rect 191104 249552 191156 249558
rect 191104 249494 191156 249500
rect 191104 249212 191156 249218
rect 191104 249154 191156 249160
rect 189460 241454 189842 241482
rect 191116 241468 191144 249154
rect 193140 243982 193168 369854
rect 193220 339040 193272 339046
rect 193220 338982 193272 338988
rect 192300 243976 192352 243982
rect 192300 243918 192352 243924
rect 193128 243976 193180 243982
rect 193128 243918 193180 243924
rect 192312 241468 192340 243918
rect 193232 241482 193260 338982
rect 193876 251122 193904 700334
rect 196624 524476 196676 524482
rect 196624 524418 196676 524424
rect 195244 334892 195296 334898
rect 195244 334834 195296 334840
rect 193864 251116 193916 251122
rect 193864 251058 193916 251064
rect 195256 243778 195284 334834
rect 196636 262886 196664 524418
rect 198648 372632 198700 372638
rect 198648 372574 198700 372580
rect 196624 262880 196676 262886
rect 196624 262822 196676 262828
rect 198660 243982 198688 372574
rect 200764 334960 200816 334966
rect 200764 334902 200816 334908
rect 200776 243982 200804 334902
rect 201512 252414 201540 702986
rect 211804 700460 211856 700466
rect 211804 700402 211856 700408
rect 207664 683188 207716 683194
rect 207664 683130 207716 683136
rect 204904 576904 204956 576910
rect 204904 576846 204956 576852
rect 203524 337204 203576 337210
rect 203524 337146 203576 337152
rect 201500 252408 201552 252414
rect 201500 252350 201552 252356
rect 203536 244254 203564 337146
rect 204916 246974 204944 576846
rect 207676 247042 207704 683130
rect 209688 336116 209740 336122
rect 209688 336058 209740 336064
rect 207664 247036 207716 247042
rect 207664 246978 207716 246984
rect 204904 246968 204956 246974
rect 204904 246910 204956 246916
rect 209700 244254 209728 336058
rect 211816 252346 211844 700402
rect 216588 337340 216640 337346
rect 216588 337282 216640 337288
rect 213184 336388 213236 336394
rect 213184 336330 213236 336336
rect 211804 252340 211856 252346
rect 211804 252282 211856 252288
rect 202328 244248 202380 244254
rect 202328 244190 202380 244196
rect 203524 244248 203576 244254
rect 203524 244190 203576 244196
rect 208676 244248 208728 244254
rect 208676 244190 208728 244196
rect 209688 244248 209740 244254
rect 209688 244190 209740 244196
rect 197360 243976 197412 243982
rect 197360 243918 197412 243924
rect 198648 243976 198700 243982
rect 198648 243918 198700 243924
rect 200764 243976 200816 243982
rect 200764 243918 200816 243924
rect 196072 243908 196124 243914
rect 196072 243850 196124 243856
rect 194876 243772 194928 243778
rect 194876 243714 194928 243720
rect 195244 243772 195296 243778
rect 195244 243714 195296 243720
rect 193232 241454 193614 241482
rect 194888 241468 194916 243714
rect 196084 241468 196112 243850
rect 197372 241468 197400 243918
rect 198648 243704 198700 243710
rect 198648 243646 198700 243652
rect 198660 241468 198688 243646
rect 201132 243500 201184 243506
rect 201132 243442 201184 243448
rect 199844 243432 199896 243438
rect 199844 243374 199896 243380
rect 199856 241468 199884 243374
rect 201144 241468 201172 243442
rect 202340 241468 202368 244190
rect 206100 244180 206152 244186
rect 206100 244122 206152 244128
rect 204904 243772 204956 243778
rect 204904 243714 204956 243720
rect 203616 243704 203668 243710
rect 203616 243646 203668 243652
rect 203628 241468 203656 243646
rect 204916 241468 204944 243714
rect 206112 241468 206140 244122
rect 207388 243908 207440 243914
rect 207388 243850 207440 243856
rect 207400 241468 207428 243850
rect 208688 241468 208716 244190
rect 213196 244186 213224 336330
rect 214564 336252 214616 336258
rect 214564 336194 214616 336200
rect 213184 244180 213236 244186
rect 213184 244122 213236 244128
rect 213644 243976 213696 243982
rect 213644 243918 213696 243924
rect 211160 243908 211212 243914
rect 211160 243850 211212 243856
rect 209872 243500 209924 243506
rect 209872 243442 209924 243448
rect 209884 241468 209912 243442
rect 211172 241468 211200 243850
rect 212448 243364 212500 243370
rect 212448 243306 212500 243312
rect 212460 241468 212488 243306
rect 213656 241468 213684 243918
rect 214576 243846 214604 336194
rect 214932 243976 214984 243982
rect 214932 243918 214984 243924
rect 214564 243840 214616 243846
rect 214564 243782 214616 243788
rect 214944 241468 214972 243918
rect 216600 241482 216628 337282
rect 218072 246158 218100 703582
rect 218808 703474 218836 703582
rect 218950 703520 219062 704960
rect 234632 703582 235028 703610
rect 218992 703474 219020 703520
rect 218808 703446 219020 703474
rect 226984 337748 227036 337754
rect 226984 337690 227036 337696
rect 225604 337680 225656 337686
rect 225604 337622 225656 337628
rect 221464 337408 221516 337414
rect 221464 337350 221516 337356
rect 220084 333464 220136 333470
rect 220084 333406 220136 333412
rect 218152 246696 218204 246702
rect 218152 246638 218204 246644
rect 218060 246152 218112 246158
rect 218060 246094 218112 246100
rect 218164 242978 218192 246638
rect 219900 244044 219952 244050
rect 219900 243986 219952 243992
rect 218704 243840 218756 243846
rect 218704 243782 218756 243788
rect 217888 242950 218192 242978
rect 217888 241482 217916 242950
rect 216154 241454 216628 241482
rect 217442 241454 217916 241482
rect 218716 241468 218744 243782
rect 219912 241468 219940 243986
rect 220096 243098 220124 333406
rect 220820 253564 220872 253570
rect 220820 253506 220872 253512
rect 220084 243092 220136 243098
rect 220084 243034 220136 243040
rect 220832 241482 220860 253506
rect 220832 241454 221214 241482
rect 221476 241058 221504 337350
rect 222844 265668 222896 265674
rect 222844 265610 222896 265616
rect 222476 244112 222528 244118
rect 222476 244054 222528 244060
rect 222488 241468 222516 244054
rect 222856 243370 222884 265610
rect 223672 244928 223724 244934
rect 223672 244870 223724 244876
rect 222844 243364 222896 243370
rect 222844 243306 222896 243312
rect 223684 241468 223712 244870
rect 224960 244044 225012 244050
rect 224960 243986 225012 243992
rect 224972 241468 225000 243986
rect 225616 243506 225644 337622
rect 226996 244186 227024 337690
rect 234528 337136 234580 337142
rect 234528 337078 234580 337084
rect 229744 336252 229796 336258
rect 229744 336194 229796 336200
rect 226984 244180 227036 244186
rect 226984 244122 227036 244128
rect 228732 244112 228784 244118
rect 228732 244054 228784 244060
rect 225604 243500 225656 243506
rect 225604 243442 225656 243448
rect 226248 243364 226300 243370
rect 226248 243306 226300 243312
rect 226260 241468 226288 243306
rect 227444 243092 227496 243098
rect 227444 243034 227496 243040
rect 227456 241468 227484 243034
rect 228744 241468 228772 244054
rect 229756 243438 229784 336194
rect 232504 273964 232556 273970
rect 232504 273906 232556 273912
rect 230480 271176 230532 271182
rect 230480 271118 230532 271124
rect 230492 267734 230520 271118
rect 230492 267706 230888 267734
rect 229928 244112 229980 244118
rect 229928 244054 229980 244060
rect 229744 243432 229796 243438
rect 229744 243374 229796 243380
rect 229940 241468 229968 244054
rect 230860 241482 230888 267706
rect 232228 243500 232280 243506
rect 232228 243442 232280 243448
rect 232240 241482 232268 243442
rect 232516 243234 232544 273906
rect 234540 244254 234568 337078
rect 234632 245206 234660 703582
rect 235000 703474 235028 703582
rect 235142 703520 235254 704960
rect 251426 703520 251538 704960
rect 267618 703520 267730 704960
rect 283810 703520 283922 704960
rect 299492 703582 299980 703610
rect 235184 703474 235212 703520
rect 235000 703446 235212 703474
rect 262864 700324 262916 700330
rect 262864 700266 262916 700272
rect 258724 590708 258776 590714
rect 258724 590650 258776 590656
rect 255964 510672 256016 510678
rect 255964 510614 256016 510620
rect 254584 375420 254636 375426
rect 254584 375362 254636 375368
rect 251824 372700 251876 372706
rect 251824 372642 251876 372648
rect 250444 369980 250496 369986
rect 250444 369922 250496 369928
rect 249064 367124 249116 367130
rect 249064 367066 249116 367072
rect 236644 337884 236696 337890
rect 236644 337826 236696 337832
rect 234620 245200 234672 245206
rect 234620 245142 234672 245148
rect 233700 244248 233752 244254
rect 233700 244190 233752 244196
rect 234528 244248 234580 244254
rect 234528 244190 234580 244196
rect 232504 243228 232556 243234
rect 232504 243170 232556 243176
rect 230860 241454 231242 241482
rect 232240 241454 232530 241482
rect 233712 241468 233740 244190
rect 236276 244180 236328 244186
rect 236276 244122 236328 244128
rect 234988 243228 235040 243234
rect 234988 243170 235040 243176
rect 235000 241468 235028 243170
rect 236288 241468 236316 244122
rect 236656 241194 236684 337826
rect 239404 337612 239456 337618
rect 239404 337554 239456 337560
rect 238760 244248 238812 244254
rect 238760 244190 238812 244196
rect 237472 244180 237524 244186
rect 237472 244122 237524 244128
rect 237484 241468 237512 244122
rect 238772 241468 238800 244190
rect 236644 241188 236696 241194
rect 236644 241130 236696 241136
rect 221464 241052 221516 241058
rect 221464 240994 221516 241000
rect 187700 240984 187752 240990
rect 187700 240926 187752 240932
rect 177028 240916 177330 240922
rect 177080 240910 177330 240916
rect 180892 240916 181102 240922
rect 177028 240858 177080 240864
rect 180944 240910 181102 240916
rect 182088 240916 182298 240922
rect 180892 240858 180944 240864
rect 182140 240910 182298 240916
rect 184664 240916 184716 240922
rect 182088 240858 182140 240864
rect 184664 240858 184716 240864
rect 40500 186448 40552 186454
rect 40500 186390 40552 186396
rect 40696 38622 40724 40052
rect 42076 39953 42104 40052
rect 42062 39944 42118 39953
rect 42062 39879 42118 39888
rect 40684 38616 40736 38622
rect 42076 38593 42104 39879
rect 40684 38558 40736 38564
rect 42062 38584 42118 38593
rect 40408 38480 40460 38486
rect 40408 38422 40460 38428
rect 39488 38412 39540 38418
rect 39488 38354 39540 38360
rect 37096 38072 37148 38078
rect 37096 38014 37148 38020
rect 19984 37188 20036 37194
rect 19984 37130 20036 37136
rect 15844 36916 15896 36922
rect 15844 36858 15896 36864
rect 14464 20664 14516 20670
rect 14464 20606 14516 20612
rect 13556 6886 13768 6914
rect 10324 6860 10376 6866
rect 10324 6802 10376 6808
rect 10322 6216 10378 6225
rect 10322 6151 10378 6160
rect 9956 4820 10008 4826
rect 9956 4762 10008 4768
rect 7656 3528 7708 3534
rect 7656 3470 7708 3476
rect 8208 3528 8260 3534
rect 8208 3470 8260 3476
rect 7668 480 7696 3470
rect 8760 3392 8812 3398
rect 8760 3334 8812 3340
rect 8772 480 8800 3334
rect 9968 480 9996 4762
rect 10336 3602 10364 6151
rect 11152 3936 11204 3942
rect 11152 3878 11204 3884
rect 10324 3596 10376 3602
rect 10324 3538 10376 3544
rect 11164 480 11192 3878
rect 12348 3596 12400 3602
rect 12348 3538 12400 3544
rect 12360 480 12388 3538
rect 13556 480 13584 6886
rect 14740 3868 14792 3874
rect 14740 3810 14792 3816
rect 14752 480 14780 3810
rect 15856 3466 15884 36858
rect 17868 36712 17920 36718
rect 17868 36654 17920 36660
rect 15936 3732 15988 3738
rect 15936 3674 15988 3680
rect 15844 3460 15896 3466
rect 15844 3402 15896 3408
rect 15948 480 15976 3674
rect 17880 3534 17908 36654
rect 19432 4072 19484 4078
rect 19432 4014 19484 4020
rect 17040 3528 17092 3534
rect 17040 3470 17092 3476
rect 17868 3528 17920 3534
rect 17868 3470 17920 3476
rect 17052 480 17080 3470
rect 18236 2916 18288 2922
rect 18236 2858 18288 2864
rect 18248 480 18276 2858
rect 19444 480 19472 4014
rect 19996 3602 20024 37130
rect 32404 37052 32456 37058
rect 32404 36994 32456 37000
rect 22008 36644 22060 36650
rect 22008 36586 22060 36592
rect 22020 6914 22048 36586
rect 25504 35556 25556 35562
rect 25504 35498 25556 35504
rect 24124 35352 24176 35358
rect 24124 35294 24176 35300
rect 21836 6886 22048 6914
rect 19984 3596 20036 3602
rect 19984 3538 20036 3544
rect 20628 3460 20680 3466
rect 20628 3402 20680 3408
rect 20640 480 20668 3402
rect 21836 480 21864 6886
rect 23020 3528 23072 3534
rect 23020 3470 23072 3476
rect 23032 480 23060 3470
rect 24136 3398 24164 35294
rect 24768 7608 24820 7614
rect 24768 7550 24820 7556
rect 24216 4004 24268 4010
rect 24216 3946 24268 3952
rect 24124 3392 24176 3398
rect 24124 3334 24176 3340
rect 24228 480 24256 3946
rect 24780 3534 24808 7550
rect 25320 3596 25372 3602
rect 25320 3538 25372 3544
rect 24768 3528 24820 3534
rect 24768 3470 24820 3476
rect 25332 480 25360 3538
rect 25516 2922 25544 35498
rect 28908 35420 28960 35426
rect 28908 35362 28960 35368
rect 28920 3466 28948 35362
rect 31668 35284 31720 35290
rect 31668 35226 31720 35232
rect 31680 6914 31708 35226
rect 31312 6886 31708 6914
rect 29000 5024 29052 5030
rect 29000 4966 29052 4972
rect 27712 3460 27764 3466
rect 27712 3402 27764 3408
rect 28908 3460 28960 3466
rect 28908 3402 28960 3408
rect 25504 2916 25556 2922
rect 25504 2858 25556 2864
rect 26516 2848 26568 2854
rect 26516 2790 26568 2796
rect 26528 480 26556 2790
rect 27724 480 27752 3402
rect 28908 3324 28960 3330
rect 28908 3266 28960 3272
rect 28920 480 28948 3266
rect 29012 2854 29040 4966
rect 30104 3664 30156 3670
rect 30104 3606 30156 3612
rect 29000 2848 29052 2854
rect 29000 2790 29052 2796
rect 30116 480 30144 3606
rect 31312 480 31340 6886
rect 32416 3670 32444 36994
rect 34428 36984 34480 36990
rect 34428 36926 34480 36932
rect 32404 3664 32456 3670
rect 32404 3606 32456 3612
rect 34440 3466 34468 36926
rect 35808 35488 35860 35494
rect 35808 35430 35860 35436
rect 35820 3466 35848 35430
rect 37108 3466 37136 38014
rect 39948 38004 40000 38010
rect 39948 37946 40000 37952
rect 38568 36848 38620 36854
rect 38568 36790 38620 36796
rect 38580 6914 38608 36790
rect 39960 6914 39988 37946
rect 40696 36582 40724 38558
rect 42062 38519 42118 38528
rect 43456 37074 43484 40052
rect 43364 37046 43484 37074
rect 43364 36922 43392 37046
rect 43352 36916 43404 36922
rect 43352 36858 43404 36864
rect 43444 36916 43496 36922
rect 43444 36858 43496 36864
rect 40684 36576 40736 36582
rect 40684 36518 40736 36524
rect 38396 6886 38608 6914
rect 39592 6886 39988 6914
rect 37188 4888 37240 4894
rect 37188 4830 37240 4836
rect 33600 3460 33652 3466
rect 33600 3402 33652 3408
rect 34428 3460 34480 3466
rect 34428 3402 34480 3408
rect 34796 3460 34848 3466
rect 34796 3402 34848 3408
rect 35808 3460 35860 3466
rect 35808 3402 35860 3408
rect 35992 3460 36044 3466
rect 35992 3402 36044 3408
rect 37096 3460 37148 3466
rect 37096 3402 37148 3408
rect 32404 3392 32456 3398
rect 32404 3334 32456 3340
rect 32416 480 32444 3334
rect 33612 480 33640 3402
rect 34808 480 34836 3402
rect 36004 480 36032 3402
rect 37200 480 37228 4830
rect 38396 480 38424 6886
rect 39592 480 39620 6886
rect 40684 4956 40736 4962
rect 40684 4898 40736 4904
rect 40696 480 40724 4898
rect 43076 4140 43128 4146
rect 43076 4082 43128 4088
rect 41880 3460 41932 3466
rect 41880 3402 41932 3408
rect 41892 480 41920 3402
rect 43088 480 43116 4082
rect 43456 3466 43484 36858
rect 44928 36786 44956 40052
rect 44916 36780 44968 36786
rect 44916 36722 44968 36728
rect 46308 32434 46336 40052
rect 46848 37936 46900 37942
rect 46848 37878 46900 37884
rect 46296 32428 46348 32434
rect 46296 32370 46348 32376
rect 46860 6914 46888 37878
rect 47780 26234 47808 40052
rect 48964 37528 49016 37534
rect 48964 37470 49016 37476
rect 46676 6886 46888 6914
rect 46952 26206 47808 26234
rect 45468 3664 45520 3670
rect 45468 3606 45520 3612
rect 43444 3460 43496 3466
rect 43444 3402 43496 3408
rect 44272 3460 44324 3466
rect 44272 3402 44324 3408
rect 44284 480 44312 3402
rect 45480 480 45508 3606
rect 46676 480 46704 6886
rect 46952 3806 46980 26206
rect 47860 6316 47912 6322
rect 47860 6258 47912 6264
rect 46940 3800 46992 3806
rect 46940 3742 46992 3748
rect 47872 480 47900 6258
rect 48976 4826 49004 37470
rect 49160 37126 49188 40052
rect 49148 37120 49200 37126
rect 49148 37062 49200 37068
rect 50632 35358 50660 40052
rect 51724 37868 51776 37874
rect 51724 37810 51776 37816
rect 50620 35352 50672 35358
rect 50620 35294 50672 35300
rect 50988 35352 51040 35358
rect 50988 35294 51040 35300
rect 48964 4820 49016 4826
rect 48964 4762 49016 4768
rect 48964 3800 49016 3806
rect 48964 3742 49016 3748
rect 48976 480 49004 3742
rect 51000 3330 51028 35294
rect 51356 6384 51408 6390
rect 51356 6326 51408 6332
rect 50160 3324 50212 3330
rect 50160 3266 50212 3272
rect 50988 3324 51040 3330
rect 50988 3266 51040 3272
rect 50172 480 50200 3266
rect 51368 480 51396 6326
rect 51736 3942 51764 37810
rect 52012 37534 52040 40052
rect 53484 37874 53512 40052
rect 53472 37868 53524 37874
rect 53472 37810 53524 37816
rect 52000 37528 52052 37534
rect 52000 37470 52052 37476
rect 54484 37324 54536 37330
rect 54484 37266 54536 37272
rect 53748 36780 53800 36786
rect 53748 36722 53800 36728
rect 51724 3936 51776 3942
rect 51724 3878 51776 3884
rect 52552 3936 52604 3942
rect 52552 3878 52604 3884
rect 52564 480 52592 3878
rect 53760 480 53788 36722
rect 54496 4078 54524 37266
rect 54864 37194 54892 40052
rect 56336 38026 56364 40052
rect 55232 37998 56364 38026
rect 54852 37188 54904 37194
rect 54852 37130 54904 37136
rect 55232 35222 55260 37998
rect 55864 37732 55916 37738
rect 55864 37674 55916 37680
rect 55220 35216 55272 35222
rect 55220 35158 55272 35164
rect 54944 6248 54996 6254
rect 54944 6190 54996 6196
rect 54484 4072 54536 4078
rect 54484 4014 54536 4020
rect 54956 480 54984 6190
rect 55876 3874 55904 37674
rect 57716 37330 57744 40052
rect 59188 37874 59216 40052
rect 60004 38276 60056 38282
rect 60004 38218 60056 38224
rect 57980 37868 58032 37874
rect 57980 37810 58032 37816
rect 59176 37868 59228 37874
rect 59176 37810 59228 37816
rect 57704 37324 57756 37330
rect 57704 37266 57756 37272
rect 57888 36576 57940 36582
rect 57888 36518 57940 36524
rect 56048 4820 56100 4826
rect 56048 4762 56100 4768
rect 55864 3868 55916 3874
rect 55864 3810 55916 3816
rect 56060 480 56088 4762
rect 57900 3330 57928 36518
rect 57992 3738 58020 37810
rect 60016 4010 60044 38218
rect 60568 36718 60596 40052
rect 61384 38140 61436 38146
rect 61384 38082 61436 38088
rect 60740 37868 60792 37874
rect 60740 37810 60792 37816
rect 60556 36712 60608 36718
rect 60556 36654 60608 36660
rect 60752 35562 60780 37810
rect 60740 35556 60792 35562
rect 60740 35498 60792 35504
rect 60004 4004 60056 4010
rect 60004 3946 60056 3952
rect 59636 3868 59688 3874
rect 59636 3810 59688 3816
rect 57980 3732 58032 3738
rect 57980 3674 58032 3680
rect 57244 3324 57296 3330
rect 57244 3266 57296 3272
rect 57888 3324 57940 3330
rect 57888 3266 57940 3272
rect 58440 3324 58492 3330
rect 58440 3266 58492 3272
rect 57256 480 57284 3266
rect 58452 480 58480 3266
rect 59648 480 59676 3810
rect 60832 3732 60884 3738
rect 60832 3674 60884 3680
rect 60844 480 60872 3674
rect 61396 3262 61424 38082
rect 62040 37874 62068 40052
rect 62028 37868 62080 37874
rect 62028 37810 62080 37816
rect 63420 37738 63448 40052
rect 63408 37732 63460 37738
rect 63408 37674 63460 37680
rect 64788 35216 64840 35222
rect 64788 35158 64840 35164
rect 61660 6588 61712 6594
rect 61660 6530 61712 6536
rect 61672 3330 61700 6530
rect 62028 6180 62080 6186
rect 62028 6122 62080 6128
rect 61660 3324 61712 3330
rect 61660 3266 61712 3272
rect 61384 3256 61436 3262
rect 61384 3198 61436 3204
rect 62040 480 62068 6122
rect 63224 4004 63276 4010
rect 63224 3946 63276 3952
rect 63236 480 63264 3946
rect 64800 3330 64828 35158
rect 64892 3534 64920 40052
rect 66272 36650 66300 40052
rect 66904 38208 66956 38214
rect 66904 38150 66956 38156
rect 66260 36644 66312 36650
rect 66260 36586 66312 36592
rect 66720 4684 66772 4690
rect 66720 4626 66772 4632
rect 64880 3528 64932 3534
rect 64880 3470 64932 3476
rect 65524 3528 65576 3534
rect 65524 3470 65576 3476
rect 64328 3324 64380 3330
rect 64328 3266 64380 3272
rect 64788 3324 64840 3330
rect 64788 3266 64840 3272
rect 64340 480 64368 3266
rect 65536 480 65564 3470
rect 66732 480 66760 4626
rect 66916 3398 66944 38150
rect 67744 26234 67772 40052
rect 69124 38282 69152 40052
rect 69112 38276 69164 38282
rect 69112 38218 69164 38224
rect 70596 37738 70624 40052
rect 69664 37732 69716 37738
rect 69664 37674 69716 37680
rect 70584 37732 70636 37738
rect 70584 37674 70636 37680
rect 68284 36712 68336 36718
rect 68284 36654 68336 36660
rect 67652 26206 67772 26234
rect 67652 7614 67680 26206
rect 67640 7608 67692 7614
rect 67640 7550 67692 7556
rect 67916 4004 67968 4010
rect 67916 3946 67968 3952
rect 66904 3392 66956 3398
rect 66904 3334 66956 3340
rect 67928 480 67956 3946
rect 68296 3534 68324 36654
rect 69676 3602 69704 37674
rect 71044 36644 71096 36650
rect 71044 36586 71096 36592
rect 70308 5364 70360 5370
rect 70308 5306 70360 5312
rect 69664 3596 69716 3602
rect 69664 3538 69716 3544
rect 68284 3528 68336 3534
rect 68284 3470 68336 3476
rect 69112 3528 69164 3534
rect 69112 3470 69164 3476
rect 69124 480 69152 3470
rect 70320 480 70348 5306
rect 71056 3534 71084 36586
rect 71976 26234 72004 40052
rect 73448 35426 73476 40052
rect 74828 38146 74856 40052
rect 74816 38140 74868 38146
rect 74816 38082 74868 38088
rect 75184 37188 75236 37194
rect 75184 37130 75236 37136
rect 73804 37120 73856 37126
rect 73804 37062 73856 37068
rect 73436 35420 73488 35426
rect 73436 35362 73488 35368
rect 71792 26206 72004 26234
rect 71792 5030 71820 26206
rect 73816 6914 73844 37062
rect 73724 6886 73844 6914
rect 72608 5432 72660 5438
rect 72608 5374 72660 5380
rect 71780 5024 71832 5030
rect 71780 4966 71832 4972
rect 71044 3528 71096 3534
rect 71044 3470 71096 3476
rect 71504 3392 71556 3398
rect 71504 3334 71556 3340
rect 71516 480 71544 3334
rect 72620 480 72648 5374
rect 73724 3942 73752 6886
rect 73804 4752 73856 4758
rect 73804 4694 73856 4700
rect 73712 3936 73764 3942
rect 73712 3878 73764 3884
rect 73816 480 73844 4694
rect 75000 3596 75052 3602
rect 75000 3538 75052 3544
rect 75012 480 75040 3538
rect 75196 3330 75224 37130
rect 76300 37058 76328 40052
rect 76288 37052 76340 37058
rect 76288 36994 76340 37000
rect 77680 35290 77708 40052
rect 79152 38214 79180 40052
rect 79140 38208 79192 38214
rect 79140 38150 79192 38156
rect 79324 38140 79376 38146
rect 79324 38082 79376 38088
rect 77944 35420 77996 35426
rect 77944 35362 77996 35368
rect 77668 35284 77720 35290
rect 77668 35226 77720 35232
rect 76196 5500 76248 5506
rect 76196 5442 76248 5448
rect 75184 3324 75236 3330
rect 75184 3266 75236 3272
rect 76208 480 76236 5442
rect 77392 3528 77444 3534
rect 77392 3470 77444 3476
rect 77404 480 77432 3470
rect 77956 3398 77984 35362
rect 79336 4146 79364 38082
rect 80532 36990 80560 40052
rect 80520 36984 80572 36990
rect 80520 36926 80572 36932
rect 82004 35494 82032 40052
rect 83384 38078 83412 40052
rect 83372 38072 83424 38078
rect 83372 38014 83424 38020
rect 82084 37052 82136 37058
rect 82084 36994 82136 37000
rect 81992 35488 82044 35494
rect 81992 35430 82044 35436
rect 82096 6914 82124 36994
rect 83464 36984 83516 36990
rect 83464 36926 83516 36932
rect 82004 6886 82124 6914
rect 79692 5296 79744 5302
rect 79692 5238 79744 5244
rect 79324 4140 79376 4146
rect 79324 4082 79376 4088
rect 77944 3392 77996 3398
rect 77944 3334 77996 3340
rect 78588 3324 78640 3330
rect 78588 3266 78640 3272
rect 78600 480 78628 3266
rect 79704 480 79732 5238
rect 82004 3874 82032 6886
rect 83280 5228 83332 5234
rect 83280 5170 83332 5176
rect 81992 3868 82044 3874
rect 81992 3810 82044 3816
rect 82084 3868 82136 3874
rect 82084 3810 82136 3816
rect 80888 3392 80940 3398
rect 80888 3334 80940 3340
rect 80900 480 80928 3334
rect 82096 480 82124 3810
rect 83292 480 83320 5170
rect 83476 3602 83504 36926
rect 84856 26234 84884 40052
rect 86236 36854 86264 40052
rect 87708 38010 87736 40052
rect 87696 38004 87748 38010
rect 87696 37946 87748 37952
rect 86224 36848 86276 36854
rect 86224 36790 86276 36796
rect 87604 35964 87656 35970
rect 87604 35906 87656 35912
rect 86224 35284 86276 35290
rect 86224 35226 86276 35232
rect 84212 26206 84884 26234
rect 84212 4894 84240 26206
rect 85212 6656 85264 6662
rect 85212 6598 85264 6604
rect 84200 4888 84252 4894
rect 84200 4830 84252 4836
rect 84476 3868 84528 3874
rect 84476 3810 84528 3816
rect 83464 3596 83516 3602
rect 83464 3538 83516 3544
rect 84488 480 84516 3810
rect 85224 3398 85252 6598
rect 85672 3936 85724 3942
rect 85672 3878 85724 3884
rect 85212 3392 85264 3398
rect 85212 3334 85264 3340
rect 85684 480 85712 3878
rect 86236 3806 86264 35226
rect 86868 5160 86920 5166
rect 86868 5102 86920 5108
rect 86224 3800 86276 3806
rect 86224 3742 86276 3748
rect 86880 480 86908 5102
rect 87616 3670 87644 35906
rect 89088 26234 89116 40052
rect 90364 38276 90416 38282
rect 90364 38218 90416 38224
rect 88352 26206 89116 26234
rect 88248 8968 88300 8974
rect 88248 8910 88300 8916
rect 87972 5024 88024 5030
rect 87972 4966 88024 4972
rect 87604 3664 87656 3670
rect 87604 3606 87656 3612
rect 87984 480 88012 4966
rect 88260 3534 88288 8910
rect 88352 4962 88380 26206
rect 88340 4956 88392 4962
rect 88340 4898 88392 4904
rect 90376 3534 90404 38218
rect 90560 36922 90588 40052
rect 91940 38146 91968 40052
rect 91928 38140 91980 38146
rect 91928 38082 91980 38088
rect 90548 36916 90600 36922
rect 90548 36858 90600 36864
rect 91744 36848 91796 36854
rect 91744 36790 91796 36796
rect 90456 5092 90508 5098
rect 90456 5034 90508 5040
rect 88248 3528 88300 3534
rect 88248 3470 88300 3476
rect 89168 3528 89220 3534
rect 89168 3470 89220 3476
rect 90364 3528 90416 3534
rect 90364 3470 90416 3476
rect 89180 480 89208 3470
rect 90468 2530 90496 5034
rect 91756 4078 91784 36790
rect 93320 26234 93348 40052
rect 94792 35970 94820 40052
rect 96172 37942 96200 40052
rect 96160 37936 96212 37942
rect 96160 37878 96212 37884
rect 95884 36916 95936 36922
rect 95884 36858 95936 36864
rect 94780 35964 94832 35970
rect 94780 35906 94832 35912
rect 92492 26206 93348 26234
rect 91744 4072 91796 4078
rect 91744 4014 91796 4020
rect 91560 3800 91612 3806
rect 91560 3742 91612 3748
rect 90376 2502 90496 2530
rect 90376 480 90404 2502
rect 91572 480 91600 3742
rect 92492 3466 92520 26206
rect 95332 7608 95384 7614
rect 95332 7550 95384 7556
rect 95148 4888 95200 4894
rect 95148 4830 95200 4836
rect 92756 4072 92808 4078
rect 92756 4014 92808 4020
rect 92480 3460 92532 3466
rect 92480 3402 92532 3408
rect 92768 480 92796 4014
rect 93952 3528 94004 3534
rect 93952 3470 94004 3476
rect 93964 480 93992 3470
rect 95160 480 95188 4830
rect 95344 3534 95372 7550
rect 95896 3738 95924 36858
rect 97644 26234 97672 40052
rect 99024 37194 99052 40052
rect 100496 38026 100524 40052
rect 99392 37998 100524 38026
rect 99012 37188 99064 37194
rect 99012 37130 99064 37136
rect 99392 35358 99420 37998
rect 100024 37936 100076 37942
rect 100024 37878 100076 37884
rect 99380 35352 99432 35358
rect 99380 35294 99432 35300
rect 96632 26206 97672 26234
rect 96632 6322 96660 26206
rect 96620 6316 96672 6322
rect 96620 6258 96672 6264
rect 97448 6316 97500 6322
rect 97448 6258 97500 6264
rect 95884 3732 95936 3738
rect 95884 3674 95936 3680
rect 95332 3528 95384 3534
rect 95332 3470 95384 3476
rect 96252 3188 96304 3194
rect 96252 3130 96304 3136
rect 96264 480 96292 3130
rect 97460 480 97488 6258
rect 98644 3596 98696 3602
rect 98644 3538 98696 3544
rect 98656 480 98684 3538
rect 99840 3392 99892 3398
rect 99840 3334 99892 3340
rect 99852 480 99880 3334
rect 100036 3194 100064 37878
rect 101876 26234 101904 40052
rect 103348 37126 103376 40052
rect 104164 38072 104216 38078
rect 104164 38014 104216 38020
rect 103336 37120 103388 37126
rect 103336 37062 103388 37068
rect 100772 26206 101904 26234
rect 100772 6390 100800 26206
rect 100760 6384 100812 6390
rect 100760 6326 100812 6332
rect 101036 6384 101088 6390
rect 101036 6326 101088 6332
rect 100024 3188 100076 3194
rect 100024 3130 100076 3136
rect 101048 480 101076 6326
rect 102232 4956 102284 4962
rect 102232 4898 102284 4904
rect 102244 480 102272 4898
rect 104176 4146 104204 38014
rect 104728 36786 104756 40052
rect 106200 38010 106228 40052
rect 107580 38010 107608 40052
rect 108304 38140 108356 38146
rect 108304 38082 108356 38088
rect 104900 38004 104952 38010
rect 104900 37946 104952 37952
rect 106188 38004 106240 38010
rect 106188 37946 106240 37952
rect 106280 38004 106332 38010
rect 106280 37946 106332 37952
rect 107568 38004 107620 38010
rect 107568 37946 107620 37952
rect 104716 36780 104768 36786
rect 104716 36722 104768 36728
rect 104532 6452 104584 6458
rect 104532 6394 104584 6400
rect 103336 4140 103388 4146
rect 103336 4082 103388 4088
rect 104164 4140 104216 4146
rect 104164 4082 104216 4088
rect 103348 480 103376 4082
rect 104544 480 104572 6394
rect 104912 6254 104940 37946
rect 104900 6248 104952 6254
rect 104900 6190 104952 6196
rect 106292 4826 106320 37946
rect 108120 6520 108172 6526
rect 108120 6462 108172 6468
rect 106280 4820 106332 4826
rect 106280 4762 106332 4768
rect 106924 3528 106976 3534
rect 106924 3470 106976 3476
rect 105728 3460 105780 3466
rect 105728 3402 105780 3408
rect 105740 480 105768 3402
rect 106936 480 106964 3470
rect 108132 480 108160 6462
rect 108316 3534 108344 38082
rect 109052 36582 109080 40052
rect 109040 36576 109092 36582
rect 109040 36518 109092 36524
rect 110432 6594 110460 40052
rect 111904 37058 111932 40052
rect 111892 37052 111944 37058
rect 111892 36994 111944 37000
rect 113284 36922 113312 40052
rect 114756 37738 114784 40052
rect 115204 38004 115256 38010
rect 115204 37946 115256 37952
rect 113824 37732 113876 37738
rect 113824 37674 113876 37680
rect 114744 37732 114796 37738
rect 114744 37674 114796 37680
rect 113272 36916 113324 36922
rect 113272 36858 113324 36864
rect 111708 29640 111760 29646
rect 111708 29582 111760 29588
rect 111720 6914 111748 29582
rect 111628 6886 111748 6914
rect 110420 6588 110472 6594
rect 110420 6530 110472 6536
rect 109316 4820 109368 4826
rect 109316 4762 109368 4768
rect 108304 3528 108356 3534
rect 108304 3470 108356 3476
rect 109328 480 109356 4762
rect 110512 3528 110564 3534
rect 110512 3470 110564 3476
rect 110524 480 110552 3470
rect 111628 480 111656 6886
rect 113836 6186 113864 37674
rect 113824 6180 113876 6186
rect 113824 6122 113876 6128
rect 115216 3670 115244 37946
rect 116136 36854 116164 40052
rect 116124 36848 116176 36854
rect 116124 36790 116176 36796
rect 117608 35222 117636 40052
rect 118988 36718 119016 40052
rect 118976 36712 119028 36718
rect 118976 36654 119028 36660
rect 119988 36576 120040 36582
rect 119988 36518 120040 36524
rect 117596 35216 117648 35222
rect 117596 35158 117648 35164
rect 117964 34536 118016 34542
rect 117964 34478 118016 34484
rect 115296 6588 115348 6594
rect 115296 6530 115348 6536
rect 114008 3664 114060 3670
rect 114008 3606 114060 3612
rect 115204 3664 115256 3670
rect 115204 3606 115256 3612
rect 112812 3256 112864 3262
rect 112812 3198 112864 3204
rect 112824 480 112852 3198
rect 114020 480 114048 3606
rect 115308 3346 115336 6530
rect 117976 4010 118004 34478
rect 120000 6914 120028 36518
rect 120460 26234 120488 40052
rect 121840 34542 121868 40052
rect 122104 37936 122156 37942
rect 122104 37878 122156 37884
rect 121828 34536 121880 34542
rect 121828 34478 121880 34484
rect 119908 6886 120028 6914
rect 120092 26206 120488 26234
rect 118792 6248 118844 6254
rect 118792 6190 118844 6196
rect 117964 4004 118016 4010
rect 117964 3946 118016 3952
rect 117596 3732 117648 3738
rect 117596 3674 117648 3680
rect 115216 3318 115336 3346
rect 115216 480 115244 3318
rect 116400 3188 116452 3194
rect 116400 3130 116452 3136
rect 116412 480 116440 3130
rect 117608 480 117636 3674
rect 118804 480 118832 6190
rect 119908 480 119936 6886
rect 120092 4690 120120 26206
rect 120080 4684 120132 4690
rect 120080 4626 120132 4632
rect 122116 3670 122144 37878
rect 123312 36650 123340 40052
rect 123300 36644 123352 36650
rect 123300 36586 123352 36592
rect 123484 36644 123536 36650
rect 123484 36586 123536 36592
rect 123496 6914 123524 36586
rect 124692 26234 124720 40052
rect 126164 35426 126192 40052
rect 126244 35964 126296 35970
rect 126244 35906 126296 35912
rect 126152 35420 126204 35426
rect 126152 35362 126204 35368
rect 123404 6886 123524 6914
rect 124232 26206 124720 26234
rect 122288 6180 122340 6186
rect 122288 6122 122340 6128
rect 121092 3664 121144 3670
rect 121092 3606 121144 3612
rect 122104 3664 122156 3670
rect 122104 3606 122156 3612
rect 121104 480 121132 3606
rect 122300 480 122328 6122
rect 123404 3262 123432 6886
rect 124232 5370 124260 26206
rect 124220 5364 124272 5370
rect 124220 5306 124272 5312
rect 123484 4140 123536 4146
rect 123484 4082 123536 4088
rect 123392 3256 123444 3262
rect 123392 3198 123444 3204
rect 123496 480 123524 4082
rect 124680 4004 124732 4010
rect 124680 3946 124732 3952
rect 124692 480 124720 3946
rect 126256 3330 126284 35906
rect 127544 26234 127572 40052
rect 129016 26234 129044 40052
rect 130396 36990 130424 40052
rect 130384 36984 130436 36990
rect 130384 36926 130436 36932
rect 131868 26234 131896 40052
rect 133248 26234 133276 40052
rect 134720 35970 134748 40052
rect 134708 35964 134760 35970
rect 134708 35906 134760 35912
rect 136100 26234 136128 40052
rect 137572 26234 137600 40052
rect 138952 35290 138980 40052
rect 138940 35284 138992 35290
rect 138940 35226 138992 35232
rect 140424 26234 140452 40052
rect 141804 26234 141832 40052
rect 143184 26234 143212 40052
rect 144656 26234 144684 40052
rect 146036 26234 146064 40052
rect 147508 38282 147536 40052
rect 147496 38276 147548 38282
rect 147496 38218 147548 38224
rect 148888 37738 148916 40052
rect 150360 37874 150388 40052
rect 151084 38276 151136 38282
rect 151084 38218 151136 38224
rect 149060 37868 149112 37874
rect 149060 37810 149112 37816
rect 150348 37868 150400 37874
rect 150348 37810 150400 37816
rect 147680 37732 147732 37738
rect 147680 37674 147732 37680
rect 148876 37732 148928 37738
rect 148876 37674 148928 37680
rect 146944 37460 146996 37466
rect 146944 37402 146996 37408
rect 126992 26206 127572 26234
rect 128372 26206 129044 26234
rect 131132 26206 131896 26234
rect 132512 26206 133276 26234
rect 135272 26206 136128 26234
rect 136652 26206 137600 26234
rect 139412 26206 140452 26234
rect 140792 26206 141832 26234
rect 142172 26206 143212 26234
rect 143552 26206 144684 26234
rect 144932 26206 146064 26234
rect 126992 5438 127020 26206
rect 126980 5432 127032 5438
rect 126980 5374 127032 5380
rect 128372 4758 128400 26206
rect 131132 5506 131160 26206
rect 132512 8974 132540 26206
rect 132500 8968 132552 8974
rect 132500 8910 132552 8916
rect 131120 5500 131172 5506
rect 131120 5442 131172 5448
rect 135272 5302 135300 26206
rect 136652 6662 136680 26206
rect 136640 6656 136692 6662
rect 136640 6598 136692 6604
rect 135260 5296 135312 5302
rect 135260 5238 135312 5244
rect 139412 5234 139440 26206
rect 139400 5228 139452 5234
rect 139400 5170 139452 5176
rect 128360 4752 128412 4758
rect 128360 4694 128412 4700
rect 140792 3874 140820 26206
rect 142172 3942 142200 26206
rect 143552 5166 143580 26206
rect 143540 5160 143592 5166
rect 143540 5102 143592 5108
rect 144932 5030 144960 26206
rect 144920 5024 144972 5030
rect 144920 4966 144972 4972
rect 146956 4078 146984 37402
rect 147692 5098 147720 37674
rect 147680 5092 147732 5098
rect 147680 5034 147732 5040
rect 146944 4072 146996 4078
rect 146944 4014 146996 4020
rect 142160 3936 142212 3942
rect 142160 3878 142212 3884
rect 140780 3868 140832 3874
rect 140780 3810 140832 3816
rect 149072 3806 149100 37810
rect 149060 3800 149112 3806
rect 149060 3742 149112 3748
rect 151096 3398 151124 38218
rect 151740 37466 151768 40052
rect 151728 37460 151780 37466
rect 151728 37402 151780 37408
rect 153212 7614 153240 40052
rect 153200 7608 153252 7614
rect 153200 7550 153252 7556
rect 154592 4894 154620 40052
rect 156064 38214 156092 40052
rect 156052 38208 156104 38214
rect 156052 38150 156104 38156
rect 157444 26234 157472 40052
rect 158916 26234 158944 40052
rect 160296 38282 160324 40052
rect 160284 38276 160336 38282
rect 160284 38218 160336 38224
rect 160744 38208 160796 38214
rect 160744 38150 160796 38156
rect 157352 26206 157472 26234
rect 158732 26206 158944 26234
rect 157352 6322 157380 26206
rect 157340 6316 157392 6322
rect 157340 6258 157392 6264
rect 154580 4888 154632 4894
rect 154580 4830 154632 4836
rect 158732 3602 158760 26206
rect 160756 6458 160784 38150
rect 161768 26234 161796 40052
rect 163148 26234 163176 40052
rect 164620 38078 164648 40052
rect 166000 38214 166028 40052
rect 165988 38208 166040 38214
rect 165988 38150 166040 38156
rect 164608 38072 164660 38078
rect 164608 38014 164660 38020
rect 164884 38072 164936 38078
rect 164884 38014 164936 38020
rect 161492 26206 161796 26234
rect 162872 26206 163176 26234
rect 160744 6452 160796 6458
rect 160744 6394 160796 6400
rect 161492 6390 161520 26206
rect 161480 6384 161532 6390
rect 161480 6326 161532 6332
rect 162872 4962 162900 26206
rect 164896 6526 164924 38014
rect 167472 26234 167500 40052
rect 168852 38146 168880 40052
rect 168840 38140 168892 38146
rect 168840 38082 168892 38088
rect 169024 38140 169076 38146
rect 169024 38082 169076 38088
rect 167012 26206 167500 26234
rect 164884 6520 164936 6526
rect 164884 6462 164936 6468
rect 162860 4956 162912 4962
rect 162860 4898 162912 4904
rect 158720 3596 158772 3602
rect 158720 3538 158772 3544
rect 167012 3466 167040 26206
rect 169036 6594 169064 38082
rect 170324 38078 170352 40052
rect 170312 38072 170364 38078
rect 170312 38014 170364 38020
rect 171704 26234 171732 40052
rect 173176 38026 173204 40052
rect 171152 26206 171732 26234
rect 172532 37998 173204 38026
rect 169024 6588 169076 6594
rect 169024 6530 169076 6536
rect 171152 4826 171180 26206
rect 171140 4820 171192 4826
rect 171140 4762 171192 4768
rect 172532 3534 172560 37998
rect 174556 37874 174584 40052
rect 175924 38072 175976 38078
rect 175924 38014 175976 38020
rect 172612 37868 172664 37874
rect 172612 37810 172664 37816
rect 174544 37868 174596 37874
rect 174544 37810 174596 37816
rect 172624 29646 172652 37810
rect 174544 37732 174596 37738
rect 174544 37674 174596 37680
rect 172612 29640 172664 29646
rect 172612 29582 172664 29588
rect 174556 3738 174584 37674
rect 175936 4146 175964 38014
rect 176028 36650 176056 40052
rect 177408 38010 177436 40052
rect 178880 38146 178908 40052
rect 178868 38140 178920 38146
rect 178868 38082 178920 38088
rect 177396 38004 177448 38010
rect 177396 37946 177448 37952
rect 178684 38004 178736 38010
rect 178684 37946 178736 37952
rect 177304 37324 177356 37330
rect 177304 37266 177356 37272
rect 176016 36644 176068 36650
rect 176016 36586 176068 36592
rect 175924 4140 175976 4146
rect 175924 4082 175976 4088
rect 174544 3732 174596 3738
rect 174544 3674 174596 3680
rect 177316 3670 177344 37266
rect 178696 4010 178724 37946
rect 180260 37738 180288 40052
rect 180248 37732 180300 37738
rect 180248 37674 180300 37680
rect 181732 37330 181760 40052
rect 181720 37324 181772 37330
rect 181720 37266 181772 37272
rect 183112 26234 183140 40052
rect 184584 36582 184612 40052
rect 185964 37942 185992 40052
rect 185952 37936 186004 37942
rect 185952 37878 186004 37884
rect 184572 36576 184624 36582
rect 184572 36518 184624 36524
rect 187436 26234 187464 40052
rect 188816 38078 188844 40052
rect 188804 38072 188856 38078
rect 188804 38014 188856 38020
rect 190288 38010 190316 40052
rect 190276 38004 190328 38010
rect 190276 37946 190328 37952
rect 191668 35894 191696 40052
rect 193048 35894 193076 40052
rect 191668 35866 191788 35894
rect 193048 35866 193168 35894
rect 182192 26206 183140 26234
rect 186332 26206 187464 26234
rect 182192 6254 182220 26206
rect 182180 6248 182232 6254
rect 182180 6190 182232 6196
rect 186332 6186 186360 26206
rect 186320 6180 186372 6186
rect 186320 6122 186372 6128
rect 178684 4004 178736 4010
rect 178684 3946 178736 3952
rect 177304 3664 177356 3670
rect 177304 3606 177356 3612
rect 172520 3528 172572 3534
rect 172520 3470 172572 3476
rect 191760 3466 191788 35866
rect 193140 3602 193168 35866
rect 193128 3596 193180 3602
rect 193128 3538 193180 3544
rect 194520 3534 194548 40052
rect 195900 38622 195928 40052
rect 195888 38616 195940 38622
rect 195888 38558 195940 38564
rect 197372 38418 197400 40052
rect 198752 38593 198780 40052
rect 200224 38962 200252 40052
rect 200212 38956 200264 38962
rect 200212 38898 200264 38904
rect 198738 38584 198794 38593
rect 198738 38519 198794 38528
rect 197360 38412 197412 38418
rect 197360 38354 197412 38360
rect 201604 38214 201632 40052
rect 201592 38208 201644 38214
rect 201592 38150 201644 38156
rect 203076 37874 203104 40052
rect 204456 38486 204484 40052
rect 204444 38480 204496 38486
rect 204444 38422 204496 38428
rect 205928 38010 205956 40052
rect 207308 38350 207336 40052
rect 207296 38344 207348 38350
rect 207296 38286 207348 38292
rect 208780 38146 208808 40052
rect 210160 38457 210188 40052
rect 210146 38448 210202 38457
rect 210146 38383 210202 38392
rect 208768 38140 208820 38146
rect 208768 38082 208820 38088
rect 205916 38004 205968 38010
rect 205916 37946 205968 37952
rect 203064 37868 203116 37874
rect 203064 37810 203116 37816
rect 211632 37806 211660 40052
rect 213012 38554 213040 40052
rect 213000 38548 213052 38554
rect 213000 38490 213052 38496
rect 211620 37800 211672 37806
rect 211620 37742 211672 37748
rect 214484 37738 214512 40052
rect 215864 38690 215892 40052
rect 215852 38684 215904 38690
rect 215852 38626 215904 38632
rect 217336 37942 217364 40052
rect 217324 37936 217376 37942
rect 217324 37878 217376 37884
rect 214472 37732 214524 37738
rect 214472 37674 214524 37680
rect 218716 37670 218744 40052
rect 220188 39098 220216 40052
rect 220176 39092 220228 39098
rect 220176 39034 220228 39040
rect 221568 38078 221596 40052
rect 223040 38894 223068 40052
rect 223028 38888 223080 38894
rect 223028 38830 223080 38836
rect 224420 38554 224448 40052
rect 225892 38826 225920 40052
rect 225880 38820 225932 38826
rect 225880 38762 225932 38768
rect 224408 38548 224460 38554
rect 224408 38490 224460 38496
rect 227272 38486 227300 40052
rect 227260 38480 227312 38486
rect 227260 38422 227312 38428
rect 228744 38418 228772 40052
rect 230124 38758 230152 40052
rect 230112 38752 230164 38758
rect 230112 38694 230164 38700
rect 231596 38690 231624 40052
rect 232976 39030 233004 40052
rect 232964 39024 233016 39030
rect 232964 38966 233016 38972
rect 231584 38684 231636 38690
rect 231584 38626 231636 38632
rect 228732 38412 228784 38418
rect 228732 38354 228784 38360
rect 234448 38282 234476 40052
rect 235828 38593 235856 40052
rect 237300 38622 237328 40052
rect 237288 38616 237340 38622
rect 235814 38584 235870 38593
rect 237288 38558 237340 38564
rect 235814 38519 235870 38528
rect 234436 38276 234488 38282
rect 234436 38218 234488 38224
rect 221556 38072 221608 38078
rect 221556 38014 221608 38020
rect 218704 37664 218756 37670
rect 218704 37606 218756 37612
rect 238680 37602 238708 40052
rect 239416 37670 239444 337554
rect 239588 337544 239640 337550
rect 239588 337486 239640 337492
rect 239496 337476 239548 337482
rect 239496 337418 239548 337424
rect 239508 38078 239536 337418
rect 239600 38554 239628 337486
rect 239680 337272 239732 337278
rect 239680 337214 239732 337220
rect 240048 337272 240100 337278
rect 240048 337214 240100 337220
rect 239588 38548 239640 38554
rect 239588 38490 239640 38496
rect 239496 38072 239548 38078
rect 239496 38014 239548 38020
rect 239692 37738 239720 337214
rect 239772 249620 239824 249626
rect 239772 249562 239824 249568
rect 239784 238921 239812 249562
rect 240060 244254 240088 337214
rect 242900 336184 242952 336190
rect 242900 336126 242952 336132
rect 247684 336184 247736 336190
rect 247684 336126 247736 336132
rect 241520 278044 241572 278050
rect 241520 277986 241572 277992
rect 240508 250708 240560 250714
rect 240508 250650 240560 250656
rect 240140 249348 240192 249354
rect 240140 249290 240192 249296
rect 240048 244248 240100 244254
rect 240048 244190 240100 244196
rect 239770 238912 239826 238921
rect 239770 238847 239826 238856
rect 240152 38486 240180 249290
rect 240416 249280 240468 249286
rect 240416 249222 240468 249228
rect 240232 242888 240284 242894
rect 240232 242830 240284 242836
rect 240140 38480 240192 38486
rect 240140 38422 240192 38428
rect 240244 38418 240272 242830
rect 240324 242684 240376 242690
rect 240324 242626 240376 242632
rect 240336 42673 240364 242626
rect 240428 138145 240456 249222
rect 240520 154057 240548 250650
rect 240692 246900 240744 246906
rect 240692 246842 240744 246848
rect 240600 246832 240652 246838
rect 240600 246774 240652 246780
rect 240612 164665 240640 246774
rect 240704 228313 240732 246842
rect 240690 228304 240746 228313
rect 240690 228239 240746 228248
rect 240598 164656 240654 164665
rect 240598 164591 240654 164600
rect 240506 154048 240562 154057
rect 240506 153983 240562 153992
rect 240414 138136 240470 138145
rect 240414 138071 240470 138080
rect 241532 85105 241560 277986
rect 241796 247852 241848 247858
rect 241796 247794 241848 247800
rect 241612 241188 241664 241194
rect 241612 241130 241664 241136
rect 241518 85096 241574 85105
rect 241518 85031 241574 85040
rect 241520 74520 241572 74526
rect 241518 74488 241520 74497
rect 241572 74488 241574 74497
rect 241518 74423 241574 74432
rect 241520 58948 241572 58954
rect 241520 58890 241572 58896
rect 241532 58585 241560 58890
rect 241518 58576 241574 58585
rect 241518 58511 241574 58520
rect 241624 47977 241652 241130
rect 241704 241052 241756 241058
rect 241704 240994 241756 241000
rect 241716 69193 241744 240994
rect 241808 101017 241836 247794
rect 241888 241120 241940 241126
rect 241888 241062 241940 241068
rect 241900 191185 241928 241062
rect 242808 234592 242860 234598
rect 242808 234534 242860 234540
rect 242820 233617 242848 234534
rect 242806 233608 242862 233617
rect 242806 233543 242862 233552
rect 242808 223576 242860 223582
rect 242808 223518 242860 223524
rect 242820 223009 242848 223518
rect 242806 223000 242862 223009
rect 242806 222935 242862 222944
rect 242808 218000 242860 218006
rect 242808 217942 242860 217948
rect 242820 217705 242848 217942
rect 242806 217696 242862 217705
rect 242806 217631 242862 217640
rect 241980 212424 242032 212430
rect 241978 212392 241980 212401
rect 242032 212392 242034 212401
rect 241978 212327 242034 212336
rect 242532 208344 242584 208350
rect 242532 208286 242584 208292
rect 242544 207097 242572 208286
rect 242530 207088 242586 207097
rect 242530 207023 242586 207032
rect 242440 202836 242492 202842
rect 242440 202778 242492 202784
rect 242452 201793 242480 202778
rect 242438 201784 242494 201793
rect 242438 201719 242494 201728
rect 242348 197328 242400 197334
rect 242348 197270 242400 197276
rect 242360 196489 242388 197270
rect 242346 196480 242402 196489
rect 242346 196415 242402 196424
rect 241886 191176 241942 191185
rect 241886 191111 241942 191120
rect 242808 186312 242860 186318
rect 242808 186254 242860 186260
rect 242820 185881 242848 186254
rect 242806 185872 242862 185881
rect 242806 185807 242862 185816
rect 242808 180804 242860 180810
rect 242808 180746 242860 180752
rect 242820 180577 242848 180746
rect 242806 180568 242862 180577
rect 242806 180503 242862 180512
rect 242806 175264 242862 175273
rect 242806 175199 242808 175208
rect 242860 175199 242862 175208
rect 242808 175170 242860 175176
rect 241888 169992 241940 169998
rect 241886 169960 241888 169969
rect 241940 169960 241942 169969
rect 241886 169895 241942 169904
rect 241888 159452 241940 159458
rect 241888 159394 241940 159400
rect 241900 159361 241928 159394
rect 241886 159352 241942 159361
rect 241886 159287 241942 159296
rect 242808 149048 242860 149054
rect 242808 148990 242860 148996
rect 242820 148753 242848 148990
rect 242806 148744 242862 148753
rect 242806 148679 242862 148688
rect 241888 143472 241940 143478
rect 241886 143440 241888 143449
rect 241940 143440 241942 143449
rect 241886 143375 241942 143384
rect 242256 128308 242308 128314
rect 242256 128250 242308 128256
rect 242268 127537 242296 128250
rect 242254 127528 242310 127537
rect 242254 127463 242310 127472
rect 241980 122596 242032 122602
rect 241980 122538 242032 122544
rect 241992 122233 242020 122538
rect 241978 122224 242034 122233
rect 241978 122159 242034 122168
rect 242808 117292 242860 117298
rect 242808 117234 242860 117240
rect 242820 116929 242848 117234
rect 242806 116920 242862 116929
rect 242806 116855 242862 116864
rect 241888 111648 241940 111654
rect 241886 111616 241888 111625
rect 241940 111616 241942 111625
rect 241886 111551 241942 111560
rect 241888 107568 241940 107574
rect 241888 107510 241940 107516
rect 241900 106321 241928 107510
rect 241886 106312 241942 106321
rect 241886 106247 241942 106256
rect 241794 101008 241850 101017
rect 241794 100943 241850 100952
rect 242808 96008 242860 96014
rect 242808 95950 242860 95956
rect 242820 95713 242848 95950
rect 242806 95704 242862 95713
rect 242806 95639 242862 95648
rect 242806 90400 242862 90409
rect 242912 90386 242940 336126
rect 243084 334824 243136 334830
rect 243084 334766 243136 334772
rect 242992 250844 243044 250850
rect 242992 250786 243044 250792
rect 242862 90358 242940 90386
rect 242806 90335 242862 90344
rect 242256 80028 242308 80034
rect 242256 79970 242308 79976
rect 242268 79801 242296 79970
rect 242254 79792 242310 79801
rect 242254 79727 242310 79736
rect 241702 69184 241758 69193
rect 241702 69119 241758 69128
rect 242808 64864 242860 64870
rect 242808 64806 242860 64812
rect 242820 63889 242848 64806
rect 242806 63880 242862 63889
rect 242806 63815 242862 63824
rect 241980 53780 242032 53786
rect 241980 53722 242032 53728
rect 241992 53281 242020 53722
rect 241978 53272 242034 53281
rect 241978 53207 242034 53216
rect 241610 47968 241666 47977
rect 241610 47903 241666 47912
rect 240322 42664 240378 42673
rect 240322 42599 240378 42608
rect 240232 38412 240284 38418
rect 240232 38354 240284 38360
rect 239680 37732 239732 37738
rect 239680 37674 239732 37680
rect 239404 37664 239456 37670
rect 239404 37606 239456 37612
rect 243004 37602 243032 250786
rect 243096 132841 243124 334766
rect 244464 333328 244516 333334
rect 244464 333270 244516 333276
rect 243452 253496 243504 253502
rect 243452 253438 243504 253444
rect 243176 252068 243228 252074
rect 243176 252010 243228 252016
rect 243082 132832 243138 132841
rect 243082 132767 243138 132776
rect 243188 74526 243216 252010
rect 243360 242820 243412 242826
rect 243360 242762 243412 242768
rect 243268 242752 243320 242758
rect 243268 242694 243320 242700
rect 243280 111654 243308 242694
rect 243372 159458 243400 242762
rect 243464 212430 243492 253438
rect 244372 242208 244424 242214
rect 244372 242150 244424 242156
rect 244280 242140 244332 242146
rect 244280 242082 244332 242088
rect 243452 212424 243504 212430
rect 243452 212366 243504 212372
rect 243360 159452 243412 159458
rect 243360 159394 243412 159400
rect 243268 111648 243320 111654
rect 243268 111590 243320 111596
rect 243176 74520 243228 74526
rect 243176 74462 243228 74468
rect 244292 38622 244320 242082
rect 244384 58954 244412 242150
rect 244476 169998 244504 333270
rect 244648 269816 244700 269822
rect 244648 269758 244700 269764
rect 244556 254652 244608 254658
rect 244556 254594 244608 254600
rect 244464 169992 244516 169998
rect 244464 169934 244516 169940
rect 244568 107574 244596 254594
rect 244660 143478 244688 269758
rect 245660 254584 245712 254590
rect 245660 254526 245712 254532
rect 244648 143472 244700 143478
rect 244648 143414 244700 143420
rect 245672 122602 245700 254526
rect 245660 122596 245712 122602
rect 245660 122538 245712 122544
rect 244556 107568 244608 107574
rect 244556 107510 244608 107516
rect 244372 58948 244424 58954
rect 244372 58890 244424 58896
rect 244280 38616 244332 38622
rect 244280 38558 244332 38564
rect 247696 38214 247724 336126
rect 249076 80034 249104 367066
rect 250456 96014 250484 369922
rect 250444 96008 250496 96014
rect 250444 95950 250496 95956
rect 249064 80028 249116 80034
rect 249064 79970 249116 79976
rect 247684 38208 247736 38214
rect 247684 38150 247736 38156
rect 251836 38146 251864 372642
rect 254596 117298 254624 375362
rect 255976 250646 256004 510614
rect 258736 260166 258764 590650
rect 261484 376780 261536 376786
rect 261484 376722 261536 376728
rect 258724 260160 258776 260166
rect 258724 260102 258776 260108
rect 255964 250640 256016 250646
rect 255964 250582 256016 250588
rect 261496 247790 261524 376722
rect 262876 264314 262904 700266
rect 267660 697610 267688 703520
rect 283852 702434 283880 703520
rect 282932 702406 283880 702434
rect 266360 697604 266412 697610
rect 266360 697546 266412 697552
rect 267648 697604 267700 697610
rect 267648 697546 267700 697552
rect 262864 264308 262916 264314
rect 262864 264250 262916 264256
rect 266372 252142 266400 697546
rect 266360 252136 266412 252142
rect 266360 252078 266412 252084
rect 261484 247784 261536 247790
rect 261484 247726 261536 247732
rect 282932 246770 282960 702406
rect 282920 246764 282972 246770
rect 282920 246706 282972 246712
rect 299492 245002 299520 703582
rect 299952 703474 299980 703582
rect 300094 703520 300206 704960
rect 316286 703520 316398 704960
rect 332478 703520 332590 704960
rect 348762 703520 348874 704960
rect 364954 703520 365066 704960
rect 381146 703520 381258 704960
rect 397430 703520 397542 704960
rect 413622 703520 413734 704960
rect 429814 703520 429926 704960
rect 446098 703520 446210 704960
rect 462290 703520 462402 704960
rect 478482 703520 478594 704960
rect 494766 703520 494878 704960
rect 510958 703520 511070 704960
rect 527150 703520 527262 704960
rect 543434 703520 543546 704960
rect 559626 703520 559738 704960
rect 575818 703520 575930 704960
rect 300136 703474 300164 703520
rect 299952 703446 300164 703474
rect 327724 700596 327776 700602
rect 327724 700538 327776 700544
rect 327736 253366 327764 700538
rect 330484 700528 330536 700534
rect 330484 700470 330536 700476
rect 327724 253360 327776 253366
rect 327724 253302 327776 253308
rect 330496 250578 330524 700470
rect 332520 700398 332548 703520
rect 333244 700664 333296 700670
rect 333244 700606 333296 700612
rect 332508 700392 332560 700398
rect 332508 700334 332560 700340
rect 333256 256018 333284 700606
rect 348804 700466 348832 703520
rect 364996 700670 365024 703520
rect 364984 700664 365036 700670
rect 364984 700606 365036 700612
rect 348792 700460 348844 700466
rect 348792 700402 348844 700408
rect 397472 700398 397500 703520
rect 334624 700392 334676 700398
rect 334624 700334 334676 700340
rect 397460 700392 397512 700398
rect 397460 700334 397512 700340
rect 333244 256012 333296 256018
rect 333244 255954 333296 255960
rect 334636 252006 334664 700334
rect 413664 700330 413692 703520
rect 429856 700602 429884 703520
rect 429844 700596 429896 700602
rect 429844 700538 429896 700544
rect 462332 700534 462360 703520
rect 478524 702434 478552 703520
rect 477512 702406 478552 702434
rect 462320 700528 462372 700534
rect 462320 700470 462372 700476
rect 413652 700324 413704 700330
rect 413652 700266 413704 700272
rect 337658 376952 337714 376961
rect 337658 376887 337714 376896
rect 337672 376786 337700 376887
rect 337660 376780 337712 376786
rect 337660 376722 337712 376728
rect 337750 376000 337806 376009
rect 337750 375935 337806 375944
rect 337764 375426 337792 375935
rect 337752 375420 337804 375426
rect 337752 375362 337804 375368
rect 337658 373824 337714 373833
rect 337658 373759 337714 373768
rect 337474 372872 337530 372881
rect 337474 372807 337530 372816
rect 337488 372706 337516 372807
rect 337476 372700 337528 372706
rect 337476 372642 337528 372648
rect 337672 372638 337700 373759
rect 337660 372632 337712 372638
rect 337660 372574 337712 372580
rect 337474 371104 337530 371113
rect 337474 371039 337530 371048
rect 337488 369918 337516 371039
rect 337750 370016 337806 370025
rect 337750 369951 337752 369960
rect 337804 369951 337806 369960
rect 337752 369922 337804 369928
rect 337476 369912 337528 369918
rect 337476 369854 337528 369860
rect 337474 368248 337530 368257
rect 337474 368183 337530 368192
rect 337488 367130 337516 368183
rect 337476 367124 337528 367130
rect 337476 367066 337528 367072
rect 337290 350024 337346 350033
rect 337290 349959 337346 349968
rect 337304 349178 337332 349959
rect 337292 349172 337344 349178
rect 337292 349114 337344 349120
rect 337382 348392 337438 348401
rect 337382 348327 337438 348336
rect 337396 338094 337424 348327
rect 337566 348120 337622 348129
rect 337566 348055 337622 348064
rect 337384 338088 337436 338094
rect 337384 338030 337436 338036
rect 334624 252000 334676 252006
rect 334624 251942 334676 251948
rect 330484 250572 330536 250578
rect 330484 250514 330536 250520
rect 299480 244996 299532 245002
rect 299480 244938 299532 244944
rect 265624 244656 265676 244662
rect 265624 244598 265676 244604
rect 262864 244588 262916 244594
rect 262864 244530 262916 244536
rect 261484 244520 261536 244526
rect 261484 244462 261536 244468
rect 258724 244452 258776 244458
rect 258724 244394 258776 244400
rect 255964 244384 256016 244390
rect 255964 244326 256016 244332
rect 254584 117292 254636 117298
rect 254584 117234 254636 117240
rect 255976 46918 256004 244326
rect 258736 86970 258764 244394
rect 261496 126954 261524 244462
rect 262876 167006 262904 244530
rect 265636 206990 265664 244598
rect 267002 244352 267058 244361
rect 267002 244287 267058 244296
rect 265624 206984 265676 206990
rect 265624 206926 265676 206932
rect 262864 167000 262916 167006
rect 262864 166942 262916 166948
rect 261484 126948 261536 126954
rect 261484 126890 261536 126896
rect 258724 86964 258776 86970
rect 258724 86906 258776 86912
rect 255964 46912 256016 46918
rect 255964 46854 256016 46860
rect 251824 38140 251876 38146
rect 251824 38082 251876 38088
rect 238668 37596 238720 37602
rect 238668 37538 238720 37544
rect 242992 37596 243044 37602
rect 242992 37538 243044 37544
rect 267016 33114 267044 244287
rect 337580 242622 337608 348055
rect 356058 338056 356114 338065
rect 356058 337991 356114 338000
rect 368478 338056 368534 338065
rect 368478 337991 368480 338000
rect 356072 337958 356100 337991
rect 368532 337991 368534 338000
rect 371238 338056 371294 338065
rect 371238 337991 371294 338000
rect 382278 338056 382334 338065
rect 382278 337991 382334 338000
rect 386602 338056 386658 338065
rect 386602 337991 386658 338000
rect 407118 338056 407174 338065
rect 407118 337991 407174 338000
rect 368480 337962 368532 337968
rect 356060 337952 356112 337958
rect 356060 337894 356112 337900
rect 363050 337784 363106 337793
rect 363050 337719 363106 337728
rect 367098 337784 367154 337793
rect 367098 337719 367154 337728
rect 356150 337648 356206 337657
rect 356150 337583 356206 337592
rect 357438 337648 357494 337657
rect 357438 337583 357494 337592
rect 358818 337648 358874 337657
rect 358818 337583 358874 337592
rect 360198 337648 360254 337657
rect 360198 337583 360254 337592
rect 362958 337648 363014 337657
rect 362958 337583 363014 337592
rect 355324 337068 355376 337074
rect 355324 337010 355376 337016
rect 337568 242616 337620 242622
rect 337568 242558 337620 242564
rect 273904 240576 273956 240582
rect 273904 240518 273956 240524
rect 272524 240508 272576 240514
rect 272524 240450 272576 240456
rect 269764 240440 269816 240446
rect 269764 240382 269816 240388
rect 268384 240372 268436 240378
rect 268384 240314 268436 240320
rect 268396 73166 268424 240314
rect 269776 113150 269804 240382
rect 272536 153202 272564 240450
rect 273916 193186 273944 240518
rect 280804 240304 280856 240310
rect 280804 240246 280856 240252
rect 279424 240236 279476 240242
rect 279424 240178 279476 240184
rect 276664 240168 276716 240174
rect 276664 240110 276716 240116
rect 273904 193180 273956 193186
rect 273904 193122 273956 193128
rect 272524 153196 272576 153202
rect 272524 153138 272576 153144
rect 269764 113144 269816 113150
rect 269764 113086 269816 113092
rect 268384 73160 268436 73166
rect 268384 73102 268436 73108
rect 267004 33108 267056 33114
rect 267004 33050 267056 33056
rect 276676 20670 276704 240110
rect 279436 100706 279464 240178
rect 280816 139398 280844 240246
rect 280804 139392 280856 139398
rect 280804 139334 280856 139340
rect 279424 100700 279476 100706
rect 279424 100642 279476 100648
rect 355336 39098 355364 337010
rect 356164 64870 356192 337583
rect 356152 64864 356204 64870
rect 356152 64806 356204 64812
rect 357452 53786 357480 337583
rect 358832 247722 358860 337583
rect 359464 337408 359516 337414
rect 359464 337350 359516 337356
rect 359476 249218 359504 337350
rect 360212 333266 360240 337583
rect 361578 337104 361634 337113
rect 361578 337039 361634 337048
rect 361592 337006 361620 337039
rect 361580 337000 361632 337006
rect 361580 336942 361632 336948
rect 360200 333260 360252 333266
rect 360200 333202 360252 333208
rect 359464 249212 359516 249218
rect 359464 249154 359516 249160
rect 358820 247716 358872 247722
rect 358820 247658 358872 247664
rect 362972 243574 363000 337583
rect 363064 243642 363092 337719
rect 364338 337648 364394 337657
rect 364338 337583 364394 337592
rect 365718 337648 365774 337657
rect 365718 337583 365774 337592
rect 364352 275330 364380 337583
rect 364340 275324 364392 275330
rect 364340 275266 364392 275272
rect 363052 243636 363104 243642
rect 363052 243578 363104 243584
rect 362960 243568 363012 243574
rect 362960 243510 363012 243516
rect 357440 53780 357492 53786
rect 357440 53722 357492 53728
rect 355324 39092 355376 39098
rect 355324 39034 355376 39040
rect 365732 38350 365760 337583
rect 367112 38962 367140 337719
rect 367190 337648 367246 337657
rect 367190 337583 367246 337592
rect 367204 253298 367232 337583
rect 371252 337210 371280 337991
rect 378138 337920 378194 337929
rect 378138 337855 378194 337864
rect 371882 337784 371938 337793
rect 371882 337719 371938 337728
rect 376850 337784 376906 337793
rect 376850 337719 376906 337728
rect 371330 337648 371386 337657
rect 371330 337583 371386 337592
rect 371240 337204 371292 337210
rect 371240 337146 371292 337152
rect 370504 337000 370556 337006
rect 369858 336968 369914 336977
rect 367744 336932 367796 336938
rect 370504 336942 370556 336948
rect 369858 336903 369914 336912
rect 367744 336874 367796 336880
rect 367192 253292 367244 253298
rect 367192 253234 367244 253240
rect 367756 223582 367784 336874
rect 369872 336870 369900 336903
rect 369860 336864 369912 336870
rect 369860 336806 369912 336812
rect 369950 336832 370006 336841
rect 369950 336767 370006 336776
rect 369964 336190 369992 336767
rect 369952 336184 370004 336190
rect 369952 336126 370004 336132
rect 367744 223576 367796 223582
rect 367744 223518 367796 223524
rect 367100 38956 367152 38962
rect 367100 38898 367152 38904
rect 370516 38593 370544 336942
rect 370502 38584 370558 38593
rect 370502 38519 370558 38528
rect 365720 38344 365772 38350
rect 365720 38286 365772 38292
rect 371344 37806 371372 337583
rect 371896 37874 371924 337719
rect 372710 337648 372766 337657
rect 372710 337583 372766 337592
rect 373998 337648 374054 337657
rect 373998 337583 374054 337592
rect 376758 337648 376814 337657
rect 376758 337583 376814 337592
rect 372724 246634 372752 337583
rect 373264 337204 373316 337210
rect 373264 337146 373316 337152
rect 372712 246628 372764 246634
rect 372712 246570 372764 246576
rect 373276 244186 373304 337146
rect 373264 244180 373316 244186
rect 373264 244122 373316 244128
rect 374012 243710 374040 337583
rect 375378 337240 375434 337249
rect 375378 337175 375434 337184
rect 375392 337074 375420 337175
rect 375470 337104 375526 337113
rect 375380 337068 375432 337074
rect 375470 337039 375526 337048
rect 375380 337010 375432 337016
rect 374000 243704 374052 243710
rect 374000 243646 374052 243652
rect 375484 38010 375512 337039
rect 376772 242554 376800 337583
rect 376864 243914 376892 337719
rect 378152 337414 378180 337855
rect 379610 337784 379666 337793
rect 379610 337719 379666 337728
rect 379518 337648 379574 337657
rect 379518 337583 379574 337592
rect 378140 337408 378192 337414
rect 378140 337350 378192 337356
rect 377404 337068 377456 337074
rect 377404 337010 377456 337016
rect 377416 244118 377444 337010
rect 377404 244112 377456 244118
rect 377404 244054 377456 244060
rect 376852 243908 376904 243914
rect 376852 243850 376904 243856
rect 379532 243778 379560 337583
rect 379624 243846 379652 337719
rect 380990 337648 381046 337657
rect 380990 337583 381046 337592
rect 380898 337376 380954 337385
rect 380898 337311 380954 337320
rect 380912 243982 380940 337311
rect 381004 264246 381032 337583
rect 382292 337346 382320 337991
rect 385684 337680 385736 337686
rect 383658 337648 383714 337657
rect 383658 337583 383714 337592
rect 385038 337648 385094 337657
rect 385684 337622 385736 337628
rect 386418 337648 386474 337657
rect 385038 337583 385094 337592
rect 382280 337340 382332 337346
rect 382280 337282 382332 337288
rect 382924 337340 382976 337346
rect 382924 337282 382976 337288
rect 382278 337240 382334 337249
rect 382278 337175 382334 337184
rect 382292 336054 382320 337175
rect 382280 336048 382332 336054
rect 382280 335990 382332 335996
rect 380992 264240 381044 264246
rect 380992 264182 381044 264188
rect 380900 243976 380952 243982
rect 380900 243918 380952 243924
rect 379612 243840 379664 243846
rect 379612 243782 379664 243788
rect 379520 243772 379572 243778
rect 379520 243714 379572 243720
rect 376760 242548 376812 242554
rect 376760 242490 376812 242496
rect 375472 38004 375524 38010
rect 375472 37946 375524 37952
rect 382936 37942 382964 337282
rect 383672 251938 383700 337583
rect 383660 251932 383712 251938
rect 383660 251874 383712 251880
rect 385052 242486 385080 337583
rect 385130 337104 385186 337113
rect 385130 337039 385186 337048
rect 385144 336258 385172 337039
rect 385132 336252 385184 336258
rect 385132 336194 385184 336200
rect 385696 244050 385724 337622
rect 386418 337583 386474 337592
rect 385684 244044 385736 244050
rect 385684 243986 385736 243992
rect 385040 242480 385092 242486
rect 385040 242422 385092 242428
rect 386432 186318 386460 337583
rect 386616 334762 386644 337991
rect 391938 337920 391994 337929
rect 391938 337855 391994 337864
rect 394698 337920 394754 337929
rect 394698 337855 394754 337864
rect 396078 337920 396134 337929
rect 396078 337855 396134 337864
rect 398838 337920 398894 337929
rect 398838 337855 398894 337864
rect 387798 337784 387854 337793
rect 387798 337719 387854 337728
rect 390558 337784 390614 337793
rect 390558 337719 390614 337728
rect 387812 337686 387840 337719
rect 390572 337686 390600 337719
rect 387800 337680 387852 337686
rect 388444 337680 388496 337686
rect 387800 337622 387852 337628
rect 387890 337648 387946 337657
rect 387064 337612 387116 337618
rect 390560 337680 390612 337686
rect 388444 337622 388496 337628
rect 389178 337648 389234 337657
rect 387890 337583 387946 337592
rect 387064 337554 387116 337560
rect 386604 334756 386656 334762
rect 386604 334698 386656 334704
rect 387076 202842 387104 337554
rect 387904 297430 387932 337583
rect 387892 297424 387944 297430
rect 387892 297366 387944 297372
rect 388456 218006 388484 337622
rect 390560 337622 390612 337628
rect 389178 337583 389180 337592
rect 389232 337583 389234 337592
rect 389180 337554 389232 337560
rect 390558 337512 390614 337521
rect 390558 337447 390614 337456
rect 390572 337346 390600 337447
rect 390560 337340 390612 337346
rect 390560 337282 390612 337288
rect 391296 337340 391348 337346
rect 391296 337282 391348 337288
rect 391204 336796 391256 336802
rect 391204 336738 391256 336744
rect 388444 218000 388496 218006
rect 388444 217942 388496 217948
rect 387064 202836 387116 202842
rect 387064 202778 387116 202784
rect 386420 186312 386472 186318
rect 386420 186254 386472 186260
rect 391216 38282 391244 336738
rect 391308 234598 391336 337282
rect 391952 337074 391980 337855
rect 394712 337822 394740 337855
rect 394700 337816 394752 337822
rect 394700 337758 394752 337764
rect 393410 337648 393466 337657
rect 393410 337583 393466 337592
rect 391940 337068 391992 337074
rect 391940 337010 391992 337016
rect 392582 336968 392638 336977
rect 392582 336903 392638 336912
rect 391296 234592 391348 234598
rect 391296 234534 391348 234540
rect 392596 39030 392624 336903
rect 393424 128314 393452 337583
rect 393870 337512 393926 337521
rect 393870 337447 393926 337456
rect 393884 336802 393912 337447
rect 396092 337142 396120 337855
rect 396170 337648 396226 337657
rect 396170 337583 396226 337592
rect 397550 337648 397606 337657
rect 397550 337583 397606 337592
rect 396080 337136 396132 337142
rect 396080 337078 396132 337084
rect 393872 336796 393924 336802
rect 393872 336738 393924 336744
rect 396184 334694 396212 337583
rect 397458 337376 397514 337385
rect 397458 337311 397460 337320
rect 397512 337311 397514 337320
rect 397460 337282 397512 337288
rect 396172 334688 396224 334694
rect 396172 334630 396224 334636
rect 393412 128308 393464 128314
rect 393412 128250 393464 128256
rect 392584 39024 392636 39030
rect 392584 38966 392636 38972
rect 397564 38894 397592 337583
rect 398852 337278 398880 337855
rect 402978 337648 403034 337657
rect 402978 337583 403034 337592
rect 405738 337648 405794 337657
rect 405738 337583 405794 337592
rect 398840 337272 398892 337278
rect 398840 337214 398892 337220
rect 400218 336832 400274 336841
rect 400218 336767 400274 336776
rect 400232 336122 400260 336767
rect 400220 336116 400272 336122
rect 400220 336058 400272 336064
rect 397552 38888 397604 38894
rect 397552 38830 397604 38836
rect 402992 38826 403020 337583
rect 405752 149054 405780 337583
rect 407132 334626 407160 337991
rect 409878 337648 409934 337657
rect 409878 337583 409934 337592
rect 412638 337648 412694 337657
rect 412638 337583 412694 337592
rect 415398 337648 415454 337657
rect 415398 337583 415454 337592
rect 417422 337648 417478 337657
rect 417422 337583 417478 337592
rect 420918 337648 420974 337657
rect 420918 337583 420974 337592
rect 424322 337648 424378 337657
rect 424322 337583 424378 337592
rect 427818 337648 427874 337657
rect 427818 337583 427874 337592
rect 430578 337648 430634 337657
rect 430578 337583 430634 337592
rect 433338 337648 433394 337657
rect 433338 337583 433394 337592
rect 440238 337648 440294 337657
rect 440238 337583 440294 337592
rect 442998 337648 443054 337657
rect 442998 337583 443054 337592
rect 407120 334620 407172 334626
rect 407120 334562 407172 334568
rect 409892 253230 409920 337583
rect 409880 253224 409932 253230
rect 409880 253166 409932 253172
rect 412652 246702 412680 337583
rect 412640 246696 412692 246702
rect 412640 246638 412692 246644
rect 415412 175234 415440 337583
rect 417436 180810 417464 337583
rect 420184 336796 420236 336802
rect 420184 336738 420236 336744
rect 420196 244934 420224 336738
rect 420184 244928 420236 244934
rect 420184 244870 420236 244876
rect 420932 242418 420960 337583
rect 422666 336832 422722 336841
rect 422666 336767 422668 336776
rect 422720 336767 422722 336776
rect 422668 336738 422720 336744
rect 420920 242412 420972 242418
rect 420920 242354 420972 242360
rect 424336 197334 424364 337583
rect 427832 208350 427860 337583
rect 427820 208344 427872 208350
rect 427820 208286 427872 208292
rect 424324 197328 424376 197334
rect 424324 197270 424376 197276
rect 417424 180804 417476 180810
rect 417424 180746 417476 180752
rect 415400 175228 415452 175234
rect 415400 175170 415452 175176
rect 405740 149048 405792 149054
rect 405740 148990 405792 148996
rect 402980 38820 403032 38826
rect 402980 38762 403032 38768
rect 430592 38758 430620 337583
rect 430580 38752 430632 38758
rect 430580 38694 430632 38700
rect 433352 38690 433380 337583
rect 434718 337104 434774 337113
rect 434718 337039 434774 337048
rect 437478 337104 437534 337113
rect 437478 337039 437534 337048
rect 434732 336938 434760 337039
rect 437492 337006 437520 337039
rect 437480 337000 437532 337006
rect 437480 336942 437532 336948
rect 434720 336932 434772 336938
rect 434720 336874 434772 336880
rect 440252 242350 440280 337583
rect 440240 242344 440292 242350
rect 440240 242286 440292 242292
rect 443012 242282 443040 337583
rect 445758 337240 445814 337249
rect 445758 337175 445760 337184
rect 445812 337175 445814 337184
rect 445760 337146 445812 337152
rect 477512 246566 477540 702406
rect 494808 700398 494836 703520
rect 480904 700392 480956 700398
rect 480904 700334 480956 700340
rect 494796 700392 494848 700398
rect 494796 700334 494848 700340
rect 479524 700324 479576 700330
rect 479524 700266 479576 700272
rect 479536 249150 479564 700266
rect 480916 251870 480944 700334
rect 486424 418192 486476 418198
rect 486424 418134 486476 418140
rect 483664 404388 483716 404394
rect 483664 404330 483716 404336
rect 482284 351960 482336 351966
rect 482284 351902 482336 351908
rect 482296 257378 482324 351902
rect 482284 257372 482336 257378
rect 482284 257314 482336 257320
rect 480904 251864 480956 251870
rect 480904 251806 480956 251812
rect 483676 250510 483704 404330
rect 485044 364404 485096 364410
rect 485044 364346 485096 364352
rect 483664 250504 483716 250510
rect 483664 250446 483716 250452
rect 479524 249144 479576 249150
rect 479524 249086 479576 249092
rect 477500 246560 477552 246566
rect 477500 246502 477552 246508
rect 485056 246430 485084 364346
rect 486436 246498 486464 418134
rect 527192 261526 527220 703520
rect 543476 702434 543504 703520
rect 542372 702406 543504 702434
rect 527180 261520 527232 261526
rect 527180 261462 527232 261468
rect 486424 246492 486476 246498
rect 486424 246434 486476 246440
rect 485044 246424 485096 246430
rect 485044 246366 485096 246372
rect 542372 246362 542400 702406
rect 559668 700330 559696 703520
rect 559656 700324 559708 700330
rect 559656 700266 559708 700272
rect 580170 697232 580226 697241
rect 580170 697167 580226 697176
rect 580184 696998 580212 697167
rect 580172 696992 580224 696998
rect 580172 696934 580224 696940
rect 580170 683904 580226 683913
rect 580170 683839 580226 683848
rect 580184 683194 580212 683839
rect 580172 683188 580224 683194
rect 580172 683130 580224 683136
rect 580172 670744 580224 670750
rect 580170 670712 580172 670721
rect 580224 670712 580226 670721
rect 580170 670647 580226 670656
rect 580170 644056 580226 644065
rect 580170 643991 580226 644000
rect 580184 643142 580212 643991
rect 580172 643136 580224 643142
rect 580172 643078 580224 643084
rect 580262 630864 580318 630873
rect 580262 630799 580318 630808
rect 580170 617536 580226 617545
rect 580170 617471 580226 617480
rect 580184 616894 580212 617471
rect 580172 616888 580224 616894
rect 580172 616830 580224 616836
rect 580170 591016 580226 591025
rect 580170 590951 580226 590960
rect 580184 590714 580212 590951
rect 580172 590708 580224 590714
rect 580172 590650 580224 590656
rect 580170 577688 580226 577697
rect 580170 577623 580226 577632
rect 580184 576910 580212 577623
rect 580172 576904 580224 576910
rect 580172 576846 580224 576852
rect 580170 564360 580226 564369
rect 580170 564295 580226 564304
rect 580184 563106 580212 564295
rect 545764 563100 545816 563106
rect 545764 563042 545816 563048
rect 580172 563100 580224 563106
rect 580172 563042 580224 563048
rect 545776 249082 545804 563042
rect 579894 537840 579950 537849
rect 579894 537775 579950 537784
rect 579908 536858 579936 537775
rect 579896 536852 579948 536858
rect 579896 536794 579948 536800
rect 580170 524512 580226 524521
rect 580170 524447 580172 524456
rect 580224 524447 580226 524456
rect 580172 524418 580224 524424
rect 580170 511320 580226 511329
rect 580170 511255 580226 511264
rect 580184 510678 580212 511255
rect 580172 510672 580224 510678
rect 580172 510614 580224 510620
rect 580170 484664 580226 484673
rect 580170 484599 580226 484608
rect 580184 484430 580212 484599
rect 580172 484424 580224 484430
rect 580172 484366 580224 484372
rect 580170 458144 580226 458153
rect 580170 458079 580226 458088
rect 580184 456822 580212 458079
rect 580172 456816 580224 456822
rect 580172 456758 580224 456764
rect 580170 418296 580226 418305
rect 580170 418231 580226 418240
rect 580184 418198 580212 418231
rect 580172 418192 580224 418198
rect 580172 418134 580224 418140
rect 580170 404968 580226 404977
rect 580170 404903 580226 404912
rect 580184 404394 580212 404903
rect 580172 404388 580224 404394
rect 580172 404330 580224 404336
rect 580170 365120 580226 365129
rect 580170 365055 580226 365064
rect 580184 364410 580212 365055
rect 580172 364404 580224 364410
rect 580172 364346 580224 364352
rect 580172 351960 580224 351966
rect 580170 351928 580172 351937
rect 580224 351928 580226 351937
rect 580170 351863 580226 351872
rect 580276 338978 580304 630799
rect 580354 471472 580410 471481
rect 580354 471407 580410 471416
rect 580264 338972 580316 338978
rect 580264 338914 580316 338920
rect 580368 338910 580396 471407
rect 580446 431624 580502 431633
rect 580446 431559 580502 431568
rect 580356 338904 580408 338910
rect 580356 338846 580408 338852
rect 580460 338842 580488 431559
rect 580538 378448 580594 378457
rect 580538 378383 580594 378392
rect 580448 338836 580500 338842
rect 580448 338778 580500 338784
rect 580552 338774 580580 378383
rect 580540 338768 580592 338774
rect 580540 338710 580592 338716
rect 580170 325272 580226 325281
rect 580170 325207 580226 325216
rect 580184 324358 580212 325207
rect 580172 324352 580224 324358
rect 580172 324294 580224 324300
rect 580170 312080 580226 312089
rect 580170 312015 580226 312024
rect 580184 311914 580212 312015
rect 580172 311908 580224 311914
rect 580172 311850 580224 311856
rect 580170 298752 580226 298761
rect 580170 298687 580226 298696
rect 580184 298178 580212 298687
rect 580172 298172 580224 298178
rect 580172 298114 580224 298120
rect 579802 272232 579858 272241
rect 579802 272167 579858 272176
rect 579816 271930 579844 272167
rect 579804 271924 579856 271930
rect 579804 271866 579856 271872
rect 580170 258904 580226 258913
rect 580170 258839 580226 258848
rect 580184 258126 580212 258839
rect 580172 258120 580224 258126
rect 580172 258062 580224 258068
rect 545764 249076 545816 249082
rect 545764 249018 545816 249024
rect 542360 246356 542412 246362
rect 542360 246298 542412 246304
rect 579802 245576 579858 245585
rect 579802 245511 579858 245520
rect 579816 244322 579844 245511
rect 579804 244316 579856 244322
rect 579804 244258 579856 244264
rect 443000 242276 443052 242282
rect 443000 242218 443052 242224
rect 580356 240984 580408 240990
rect 580356 240926 580408 240932
rect 580264 240848 580316 240854
rect 580264 240790 580316 240796
rect 579804 240780 579856 240786
rect 579804 240722 579856 240728
rect 579816 232393 579844 240722
rect 579802 232384 579858 232393
rect 579802 232319 579858 232328
rect 579896 206984 579948 206990
rect 579896 206926 579948 206932
rect 579908 205737 579936 206926
rect 579894 205728 579950 205737
rect 579894 205663 579950 205672
rect 580172 193180 580224 193186
rect 580172 193122 580224 193128
rect 580184 192545 580212 193122
rect 580170 192536 580226 192545
rect 580170 192471 580226 192480
rect 580172 167000 580224 167006
rect 580172 166942 580224 166948
rect 580184 165889 580212 166942
rect 580170 165880 580226 165889
rect 580170 165815 580226 165824
rect 579804 153196 579856 153202
rect 579804 153138 579856 153144
rect 579816 152697 579844 153138
rect 579802 152688 579858 152697
rect 579802 152623 579858 152632
rect 580172 139392 580224 139398
rect 580170 139360 580172 139369
rect 580224 139360 580226 139369
rect 580170 139295 580226 139304
rect 580172 126948 580224 126954
rect 580172 126890 580224 126896
rect 580184 126041 580212 126890
rect 580170 126032 580226 126041
rect 580170 125967 580226 125976
rect 580172 113144 580224 113150
rect 580172 113086 580224 113092
rect 580184 112849 580212 113086
rect 580170 112840 580226 112849
rect 580170 112775 580226 112784
rect 580172 100700 580224 100706
rect 580172 100642 580224 100648
rect 580184 99521 580212 100642
rect 580170 99512 580226 99521
rect 580170 99447 580226 99456
rect 580172 86964 580224 86970
rect 580172 86906 580224 86912
rect 580184 86193 580212 86906
rect 580170 86184 580226 86193
rect 580170 86119 580226 86128
rect 579988 73160 580040 73166
rect 579988 73102 580040 73108
rect 580000 73001 580028 73102
rect 579986 72992 580042 73001
rect 579986 72927 580042 72936
rect 580276 59673 580304 240790
rect 580368 179217 580396 240926
rect 580448 240916 580500 240922
rect 580448 240858 580500 240864
rect 580460 219065 580488 240858
rect 580446 219056 580502 219065
rect 580446 218991 580502 219000
rect 580354 179208 580410 179217
rect 580354 179143 580410 179152
rect 580262 59664 580318 59673
rect 580262 59599 580318 59608
rect 580172 46912 580224 46918
rect 580172 46854 580224 46860
rect 580184 46345 580212 46854
rect 580170 46336 580226 46345
rect 580170 46271 580226 46280
rect 580264 39364 580316 39370
rect 580264 39306 580316 39312
rect 433340 38684 433392 38690
rect 433340 38626 433392 38632
rect 391204 38276 391256 38282
rect 391204 38218 391256 38224
rect 382924 37936 382976 37942
rect 382924 37878 382976 37884
rect 371884 37868 371936 37874
rect 371884 37810 371936 37816
rect 371332 37800 371384 37806
rect 371332 37742 371384 37748
rect 580170 33144 580226 33153
rect 580170 33079 580172 33088
rect 580224 33079 580226 33088
rect 580172 33050 580224 33056
rect 276664 20664 276716 20670
rect 276664 20606 276716 20612
rect 580172 20664 580224 20670
rect 580172 20606 580224 20612
rect 580184 19825 580212 20606
rect 580170 19816 580226 19825
rect 580170 19751 580226 19760
rect 580276 6633 580304 39306
rect 580262 6624 580318 6633
rect 580262 6559 580318 6568
rect 582196 3596 582248 3602
rect 582196 3538 582248 3544
rect 194508 3528 194560 3534
rect 194508 3470 194560 3476
rect 167000 3460 167052 3466
rect 167000 3402 167052 3408
rect 191748 3460 191800 3466
rect 191748 3402 191800 3408
rect 581000 3460 581052 3466
rect 581000 3402 581052 3408
rect 151084 3392 151136 3398
rect 151084 3334 151136 3340
rect 126244 3324 126296 3330
rect 126244 3266 126296 3272
rect 581012 480 581040 3402
rect 582208 480 582236 3538
rect 583392 3528 583444 3534
rect 583392 3470 583444 3476
rect 583404 480 583432 3470
rect 542 -960 654 480
rect 1646 -960 1758 480
rect 2842 -960 2954 480
rect 4038 -960 4150 480
rect 5234 -960 5346 480
rect 6430 -960 6542 480
rect 7626 -960 7738 480
rect 8730 -960 8842 480
rect 9926 -960 10038 480
rect 11122 -960 11234 480
rect 12318 -960 12430 480
rect 13514 -960 13626 480
rect 14710 -960 14822 480
rect 15906 -960 16018 480
rect 17010 -960 17122 480
rect 18206 -960 18318 480
rect 19402 -960 19514 480
rect 20598 -960 20710 480
rect 21794 -960 21906 480
rect 22990 -960 23102 480
rect 24186 -960 24298 480
rect 25290 -960 25402 480
rect 26486 -960 26598 480
rect 27682 -960 27794 480
rect 28878 -960 28990 480
rect 30074 -960 30186 480
rect 31270 -960 31382 480
rect 32374 -960 32486 480
rect 33570 -960 33682 480
rect 34766 -960 34878 480
rect 35962 -960 36074 480
rect 37158 -960 37270 480
rect 38354 -960 38466 480
rect 39550 -960 39662 480
rect 40654 -960 40766 480
rect 41850 -960 41962 480
rect 43046 -960 43158 480
rect 44242 -960 44354 480
rect 45438 -960 45550 480
rect 46634 -960 46746 480
rect 47830 -960 47942 480
rect 48934 -960 49046 480
rect 50130 -960 50242 480
rect 51326 -960 51438 480
rect 52522 -960 52634 480
rect 53718 -960 53830 480
rect 54914 -960 55026 480
rect 56018 -960 56130 480
rect 57214 -960 57326 480
rect 58410 -960 58522 480
rect 59606 -960 59718 480
rect 60802 -960 60914 480
rect 61998 -960 62110 480
rect 63194 -960 63306 480
rect 64298 -960 64410 480
rect 65494 -960 65606 480
rect 66690 -960 66802 480
rect 67886 -960 67998 480
rect 69082 -960 69194 480
rect 70278 -960 70390 480
rect 71474 -960 71586 480
rect 72578 -960 72690 480
rect 73774 -960 73886 480
rect 74970 -960 75082 480
rect 76166 -960 76278 480
rect 77362 -960 77474 480
rect 78558 -960 78670 480
rect 79662 -960 79774 480
rect 80858 -960 80970 480
rect 82054 -960 82166 480
rect 83250 -960 83362 480
rect 84446 -960 84558 480
rect 85642 -960 85754 480
rect 86838 -960 86950 480
rect 87942 -960 88054 480
rect 89138 -960 89250 480
rect 90334 -960 90446 480
rect 91530 -960 91642 480
rect 92726 -960 92838 480
rect 93922 -960 94034 480
rect 95118 -960 95230 480
rect 96222 -960 96334 480
rect 97418 -960 97530 480
rect 98614 -960 98726 480
rect 99810 -960 99922 480
rect 101006 -960 101118 480
rect 102202 -960 102314 480
rect 103306 -960 103418 480
rect 104502 -960 104614 480
rect 105698 -960 105810 480
rect 106894 -960 107006 480
rect 108090 -960 108202 480
rect 109286 -960 109398 480
rect 110482 -960 110594 480
rect 111586 -960 111698 480
rect 112782 -960 112894 480
rect 113978 -960 114090 480
rect 115174 -960 115286 480
rect 116370 -960 116482 480
rect 117566 -960 117678 480
rect 118762 -960 118874 480
rect 119866 -960 119978 480
rect 121062 -960 121174 480
rect 122258 -960 122370 480
rect 123454 -960 123566 480
rect 124650 -960 124762 480
rect 125846 -960 125958 480
rect 126950 -960 127062 480
rect 128146 -960 128258 480
rect 129342 -960 129454 480
rect 130538 -960 130650 480
rect 131734 -960 131846 480
rect 132930 -960 133042 480
rect 134126 -960 134238 480
rect 135230 -960 135342 480
rect 136426 -960 136538 480
rect 137622 -960 137734 480
rect 138818 -960 138930 480
rect 140014 -960 140126 480
rect 141210 -960 141322 480
rect 142406 -960 142518 480
rect 143510 -960 143622 480
rect 144706 -960 144818 480
rect 145902 -960 146014 480
rect 147098 -960 147210 480
rect 148294 -960 148406 480
rect 149490 -960 149602 480
rect 150594 -960 150706 480
rect 151790 -960 151902 480
rect 152986 -960 153098 480
rect 154182 -960 154294 480
rect 155378 -960 155490 480
rect 156574 -960 156686 480
rect 157770 -960 157882 480
rect 158874 -960 158986 480
rect 160070 -960 160182 480
rect 161266 -960 161378 480
rect 162462 -960 162574 480
rect 163658 -960 163770 480
rect 164854 -960 164966 480
rect 166050 -960 166162 480
rect 167154 -960 167266 480
rect 168350 -960 168462 480
rect 169546 -960 169658 480
rect 170742 -960 170854 480
rect 171938 -960 172050 480
rect 173134 -960 173246 480
rect 174238 -960 174350 480
rect 175434 -960 175546 480
rect 176630 -960 176742 480
rect 177826 -960 177938 480
rect 179022 -960 179134 480
rect 180218 -960 180330 480
rect 181414 -960 181526 480
rect 182518 -960 182630 480
rect 183714 -960 183826 480
rect 184910 -960 185022 480
rect 186106 -960 186218 480
rect 187302 -960 187414 480
rect 188498 -960 188610 480
rect 189694 -960 189806 480
rect 190798 -960 190910 480
rect 191994 -960 192106 480
rect 193190 -960 193302 480
rect 194386 -960 194498 480
rect 195582 -960 195694 480
rect 196778 -960 196890 480
rect 197882 -960 197994 480
rect 199078 -960 199190 480
rect 200274 -960 200386 480
rect 201470 -960 201582 480
rect 202666 -960 202778 480
rect 203862 -960 203974 480
rect 205058 -960 205170 480
rect 206162 -960 206274 480
rect 207358 -960 207470 480
rect 208554 -960 208666 480
rect 209750 -960 209862 480
rect 210946 -960 211058 480
rect 212142 -960 212254 480
rect 213338 -960 213450 480
rect 214442 -960 214554 480
rect 215638 -960 215750 480
rect 216834 -960 216946 480
rect 218030 -960 218142 480
rect 219226 -960 219338 480
rect 220422 -960 220534 480
rect 221526 -960 221638 480
rect 222722 -960 222834 480
rect 223918 -960 224030 480
rect 225114 -960 225226 480
rect 226310 -960 226422 480
rect 227506 -960 227618 480
rect 228702 -960 228814 480
rect 229806 -960 229918 480
rect 231002 -960 231114 480
rect 232198 -960 232310 480
rect 233394 -960 233506 480
rect 234590 -960 234702 480
rect 235786 -960 235898 480
rect 236982 -960 237094 480
rect 238086 -960 238198 480
rect 239282 -960 239394 480
rect 240478 -960 240590 480
rect 241674 -960 241786 480
rect 242870 -960 242982 480
rect 244066 -960 244178 480
rect 245170 -960 245282 480
rect 246366 -960 246478 480
rect 247562 -960 247674 480
rect 248758 -960 248870 480
rect 249954 -960 250066 480
rect 251150 -960 251262 480
rect 252346 -960 252458 480
rect 253450 -960 253562 480
rect 254646 -960 254758 480
rect 255842 -960 255954 480
rect 257038 -960 257150 480
rect 258234 -960 258346 480
rect 259430 -960 259542 480
rect 260626 -960 260738 480
rect 261730 -960 261842 480
rect 262926 -960 263038 480
rect 264122 -960 264234 480
rect 265318 -960 265430 480
rect 266514 -960 266626 480
rect 267710 -960 267822 480
rect 268814 -960 268926 480
rect 270010 -960 270122 480
rect 271206 -960 271318 480
rect 272402 -960 272514 480
rect 273598 -960 273710 480
rect 274794 -960 274906 480
rect 275990 -960 276102 480
rect 277094 -960 277206 480
rect 278290 -960 278402 480
rect 279486 -960 279598 480
rect 280682 -960 280794 480
rect 281878 -960 281990 480
rect 283074 -960 283186 480
rect 284270 -960 284382 480
rect 285374 -960 285486 480
rect 286570 -960 286682 480
rect 287766 -960 287878 480
rect 288962 -960 289074 480
rect 290158 -960 290270 480
rect 291354 -960 291466 480
rect 292550 -960 292662 480
rect 293654 -960 293766 480
rect 294850 -960 294962 480
rect 296046 -960 296158 480
rect 297242 -960 297354 480
rect 298438 -960 298550 480
rect 299634 -960 299746 480
rect 300738 -960 300850 480
rect 301934 -960 302046 480
rect 303130 -960 303242 480
rect 304326 -960 304438 480
rect 305522 -960 305634 480
rect 306718 -960 306830 480
rect 307914 -960 308026 480
rect 309018 -960 309130 480
rect 310214 -960 310326 480
rect 311410 -960 311522 480
rect 312606 -960 312718 480
rect 313802 -960 313914 480
rect 314998 -960 315110 480
rect 316194 -960 316306 480
rect 317298 -960 317410 480
rect 318494 -960 318606 480
rect 319690 -960 319802 480
rect 320886 -960 320998 480
rect 322082 -960 322194 480
rect 323278 -960 323390 480
rect 324382 -960 324494 480
rect 325578 -960 325690 480
rect 326774 -960 326886 480
rect 327970 -960 328082 480
rect 329166 -960 329278 480
rect 330362 -960 330474 480
rect 331558 -960 331670 480
rect 332662 -960 332774 480
rect 333858 -960 333970 480
rect 335054 -960 335166 480
rect 336250 -960 336362 480
rect 337446 -960 337558 480
rect 338642 -960 338754 480
rect 339838 -960 339950 480
rect 340942 -960 341054 480
rect 342138 -960 342250 480
rect 343334 -960 343446 480
rect 344530 -960 344642 480
rect 345726 -960 345838 480
rect 346922 -960 347034 480
rect 348026 -960 348138 480
rect 349222 -960 349334 480
rect 350418 -960 350530 480
rect 351614 -960 351726 480
rect 352810 -960 352922 480
rect 354006 -960 354118 480
rect 355202 -960 355314 480
rect 356306 -960 356418 480
rect 357502 -960 357614 480
rect 358698 -960 358810 480
rect 359894 -960 360006 480
rect 361090 -960 361202 480
rect 362286 -960 362398 480
rect 363482 -960 363594 480
rect 364586 -960 364698 480
rect 365782 -960 365894 480
rect 366978 -960 367090 480
rect 368174 -960 368286 480
rect 369370 -960 369482 480
rect 370566 -960 370678 480
rect 371670 -960 371782 480
rect 372866 -960 372978 480
rect 374062 -960 374174 480
rect 375258 -960 375370 480
rect 376454 -960 376566 480
rect 377650 -960 377762 480
rect 378846 -960 378958 480
rect 379950 -960 380062 480
rect 381146 -960 381258 480
rect 382342 -960 382454 480
rect 383538 -960 383650 480
rect 384734 -960 384846 480
rect 385930 -960 386042 480
rect 387126 -960 387238 480
rect 388230 -960 388342 480
rect 389426 -960 389538 480
rect 390622 -960 390734 480
rect 391818 -960 391930 480
rect 393014 -960 393126 480
rect 394210 -960 394322 480
rect 395314 -960 395426 480
rect 396510 -960 396622 480
rect 397706 -960 397818 480
rect 398902 -960 399014 480
rect 400098 -960 400210 480
rect 401294 -960 401406 480
rect 402490 -960 402602 480
rect 403594 -960 403706 480
rect 404790 -960 404902 480
rect 405986 -960 406098 480
rect 407182 -960 407294 480
rect 408378 -960 408490 480
rect 409574 -960 409686 480
rect 410770 -960 410882 480
rect 411874 -960 411986 480
rect 413070 -960 413182 480
rect 414266 -960 414378 480
rect 415462 -960 415574 480
rect 416658 -960 416770 480
rect 417854 -960 417966 480
rect 418958 -960 419070 480
rect 420154 -960 420266 480
rect 421350 -960 421462 480
rect 422546 -960 422658 480
rect 423742 -960 423854 480
rect 424938 -960 425050 480
rect 426134 -960 426246 480
rect 427238 -960 427350 480
rect 428434 -960 428546 480
rect 429630 -960 429742 480
rect 430826 -960 430938 480
rect 432022 -960 432134 480
rect 433218 -960 433330 480
rect 434414 -960 434526 480
rect 435518 -960 435630 480
rect 436714 -960 436826 480
rect 437910 -960 438022 480
rect 439106 -960 439218 480
rect 440302 -960 440414 480
rect 441498 -960 441610 480
rect 442602 -960 442714 480
rect 443798 -960 443910 480
rect 444994 -960 445106 480
rect 446190 -960 446302 480
rect 447386 -960 447498 480
rect 448582 -960 448694 480
rect 449778 -960 449890 480
rect 450882 -960 450994 480
rect 452078 -960 452190 480
rect 453274 -960 453386 480
rect 454470 -960 454582 480
rect 455666 -960 455778 480
rect 456862 -960 456974 480
rect 458058 -960 458170 480
rect 459162 -960 459274 480
rect 460358 -960 460470 480
rect 461554 -960 461666 480
rect 462750 -960 462862 480
rect 463946 -960 464058 480
rect 465142 -960 465254 480
rect 466246 -960 466358 480
rect 467442 -960 467554 480
rect 468638 -960 468750 480
rect 469834 -960 469946 480
rect 471030 -960 471142 480
rect 472226 -960 472338 480
rect 473422 -960 473534 480
rect 474526 -960 474638 480
rect 475722 -960 475834 480
rect 476918 -960 477030 480
rect 478114 -960 478226 480
rect 479310 -960 479422 480
rect 480506 -960 480618 480
rect 481702 -960 481814 480
rect 482806 -960 482918 480
rect 484002 -960 484114 480
rect 485198 -960 485310 480
rect 486394 -960 486506 480
rect 487590 -960 487702 480
rect 488786 -960 488898 480
rect 489890 -960 490002 480
rect 491086 -960 491198 480
rect 492282 -960 492394 480
rect 493478 -960 493590 480
rect 494674 -960 494786 480
rect 495870 -960 495982 480
rect 497066 -960 497178 480
rect 498170 -960 498282 480
rect 499366 -960 499478 480
rect 500562 -960 500674 480
rect 501758 -960 501870 480
rect 502954 -960 503066 480
rect 504150 -960 504262 480
rect 505346 -960 505458 480
rect 506450 -960 506562 480
rect 507646 -960 507758 480
rect 508842 -960 508954 480
rect 510038 -960 510150 480
rect 511234 -960 511346 480
rect 512430 -960 512542 480
rect 513534 -960 513646 480
rect 514730 -960 514842 480
rect 515926 -960 516038 480
rect 517122 -960 517234 480
rect 518318 -960 518430 480
rect 519514 -960 519626 480
rect 520710 -960 520822 480
rect 521814 -960 521926 480
rect 523010 -960 523122 480
rect 524206 -960 524318 480
rect 525402 -960 525514 480
rect 526598 -960 526710 480
rect 527794 -960 527906 480
rect 528990 -960 529102 480
rect 530094 -960 530206 480
rect 531290 -960 531402 480
rect 532486 -960 532598 480
rect 533682 -960 533794 480
rect 534878 -960 534990 480
rect 536074 -960 536186 480
rect 537178 -960 537290 480
rect 538374 -960 538486 480
rect 539570 -960 539682 480
rect 540766 -960 540878 480
rect 541962 -960 542074 480
rect 543158 -960 543270 480
rect 544354 -960 544466 480
rect 545458 -960 545570 480
rect 546654 -960 546766 480
rect 547850 -960 547962 480
rect 549046 -960 549158 480
rect 550242 -960 550354 480
rect 551438 -960 551550 480
rect 552634 -960 552746 480
rect 553738 -960 553850 480
rect 554934 -960 555046 480
rect 556130 -960 556242 480
rect 557326 -960 557438 480
rect 558522 -960 558634 480
rect 559718 -960 559830 480
rect 560822 -960 560934 480
rect 562018 -960 562130 480
rect 563214 -960 563326 480
rect 564410 -960 564522 480
rect 565606 -960 565718 480
rect 566802 -960 566914 480
rect 567998 -960 568110 480
rect 569102 -960 569214 480
rect 570298 -960 570410 480
rect 571494 -960 571606 480
rect 572690 -960 572802 480
rect 573886 -960 573998 480
rect 575082 -960 575194 480
rect 576278 -960 576390 480
rect 577382 -960 577494 480
rect 578578 -960 578690 480
rect 579774 -960 579886 480
rect 580970 -960 581082 480
rect 582166 -960 582278 480
rect 583362 -960 583474 480
<< via2 >>
rect 2778 684256 2834 684312
rect 3422 671200 3478 671256
rect 3330 606056 3386 606112
rect 3330 579944 3386 580000
rect 3330 553832 3386 553888
rect 3330 527856 3386 527912
rect 3330 514820 3386 514856
rect 3330 514800 3332 514820
rect 3332 514800 3384 514820
rect 3384 514800 3386 514820
rect 2870 501744 2926 501800
rect 3330 475632 3386 475688
rect 3330 462576 3386 462632
rect 3330 449520 3386 449576
rect 3146 423544 3202 423600
rect 3330 397468 3332 397488
rect 3332 397468 3384 397488
rect 3384 397468 3386 397488
rect 3330 397432 3386 397468
rect 3330 371320 3386 371376
rect 3054 345344 3110 345400
rect 3514 658144 3570 658200
rect 3514 632068 3516 632088
rect 3516 632068 3568 632088
rect 3568 632068 3570 632088
rect 3514 632032 3570 632068
rect 3514 619112 3570 619168
rect 3606 566888 3662 566944
rect 3698 410488 3754 410544
rect 3422 319232 3478 319288
rect 3422 306176 3478 306232
rect 3422 293120 3478 293176
rect 3054 267144 3110 267200
rect 3422 254088 3478 254144
rect 3790 358400 3846 358456
rect 3422 241032 3478 241088
rect 3330 214920 3386 214976
rect 3422 201864 3478 201920
rect 3422 188808 3478 188864
rect 3238 162832 3294 162888
rect 3422 149776 3478 149832
rect 3238 136720 3294 136776
rect 3422 110608 3478 110664
rect 3422 97552 3478 97608
rect 3146 84632 3202 84688
rect 3422 71576 3478 71632
rect 3054 58520 3110 58576
rect 3422 45500 3424 45520
rect 3424 45500 3476 45520
rect 3476 45500 3478 45520
rect 3422 45464 3478 45500
rect 2778 32408 2834 32464
rect 3422 19352 3478 19408
rect 3422 6432 3478 6488
rect 38474 376896 38530 376952
rect 37922 375944 37978 376000
rect 37830 348064 37886 348120
rect 36634 213016 36690 213072
rect 36726 199824 36782 199880
rect 36818 164872 36874 164928
rect 36910 156032 36966 156088
rect 37094 234912 37150 234968
rect 37186 226208 37242 226264
rect 37370 186768 37426 186824
rect 37002 142976 37058 143032
rect 37830 221720 37886 221776
rect 37738 116592 37794 116648
rect 37646 107888 37702 107944
rect 38106 373768 38162 373824
rect 38290 372816 38346 372872
rect 38382 349968 38438 350024
rect 38014 217368 38070 217424
rect 38014 195472 38070 195528
rect 38014 191120 38070 191176
rect 38014 177964 38016 177984
rect 38016 177964 38068 177984
rect 38068 177964 38070 177984
rect 38014 177928 38070 177964
rect 38014 173576 38070 173632
rect 38014 169224 38070 169280
rect 38014 160384 38070 160440
rect 38014 151716 38016 151736
rect 38016 151716 38068 151736
rect 38068 151716 38070 151736
rect 38014 151680 38070 151716
rect 38014 147328 38070 147384
rect 38014 138488 38070 138544
rect 38106 134136 38162 134192
rect 38014 129784 38070 129840
rect 38014 125432 38070 125488
rect 37922 120944 37978 121000
rect 38014 112240 38070 112296
rect 38014 94696 38070 94752
rect 38014 90344 38070 90400
rect 38014 77152 38070 77208
rect 38014 68448 38070 68504
rect 38290 99048 38346 99104
rect 38198 64096 38254 64152
rect 38014 59608 38070 59664
rect 38014 55256 38070 55312
rect 37830 50904 37886 50960
rect 38014 46552 38070 46608
rect 38014 42200 38070 42256
rect 38842 371048 38898 371104
rect 38658 369960 38714 370016
rect 38566 348336 38622 348392
rect 38750 368192 38806 368248
rect 38658 103536 38714 103592
rect 38566 85992 38622 86048
rect 39210 230560 39266 230616
rect 39118 208664 39174 208720
rect 39026 204312 39082 204368
rect 38934 182280 38990 182336
rect 38842 81504 38898 81560
rect 38750 72800 38806 72856
rect 39946 239808 40002 239864
rect 41786 244296 41842 244352
rect 56506 337884 56562 337920
rect 56506 337864 56508 337884
rect 56508 337864 56560 337884
rect 56560 337864 56562 337884
rect 68926 337728 68982 337784
rect 70582 337728 70638 337784
rect 59266 337592 59322 337648
rect 62026 337592 62082 337648
rect 63406 337592 63462 337648
rect 64970 337592 65026 337648
rect 66350 337592 66406 337648
rect 67638 337592 67694 337648
rect 57886 337456 57942 337512
rect 59450 337320 59506 337376
rect 59358 337204 59414 337240
rect 59358 337184 59360 337204
rect 59360 337184 59412 337204
rect 59412 337184 59414 337204
rect 64786 337456 64842 337512
rect 70490 337592 70546 337648
rect 69110 337320 69166 337376
rect 72974 337456 73030 337512
rect 74354 337728 74410 337784
rect 74446 337592 74502 337648
rect 74906 337592 74962 337648
rect 76286 338000 76342 338056
rect 78586 337864 78642 337920
rect 77206 337728 77262 337784
rect 78494 337592 78550 337648
rect 77206 336776 77262 336832
rect 79966 337592 80022 337648
rect 81070 337592 81126 337648
rect 81254 336776 81310 336832
rect 91006 338000 91062 338056
rect 83554 337728 83610 337784
rect 88062 337728 88118 337784
rect 82726 337592 82782 337648
rect 82910 337592 82966 337648
rect 83002 336912 83058 336968
rect 85302 337592 85358 337648
rect 86406 337592 86462 337648
rect 88154 337592 88210 337648
rect 88430 337592 88486 337648
rect 90638 337592 90694 337648
rect 91190 337592 91246 337648
rect 99286 337864 99342 337920
rect 92386 337728 92442 337784
rect 93582 337728 93638 337784
rect 95146 337728 95202 337784
rect 97998 337728 98054 337784
rect 92478 337592 92534 337648
rect 96342 337592 96398 337648
rect 97906 337592 97962 337648
rect 96526 336776 96582 336832
rect 100758 337592 100814 337648
rect 106186 337592 106242 337648
rect 107658 337592 107714 337648
rect 111706 337592 111762 337648
rect 113178 337592 113234 337648
rect 118606 337592 118662 337648
rect 121366 337592 121422 337648
rect 122838 337592 122894 337648
rect 126886 337592 126942 337648
rect 99286 336776 99342 336832
rect 104806 336776 104862 336832
rect 117226 337184 117282 337240
rect 131026 338000 131082 338056
rect 129646 337592 129702 337648
rect 132590 337592 132646 337648
rect 135258 337592 135314 337648
rect 139306 337592 139362 337648
rect 142158 337728 142214 337784
rect 142066 337592 142122 337648
rect 146206 337592 146262 337648
rect 184846 242936 184902 242992
rect 42062 39888 42118 39944
rect 10322 6160 10378 6216
rect 42062 38528 42118 38584
rect 198738 38528 198794 38584
rect 210146 38392 210202 38448
rect 235814 38528 235870 38584
rect 239770 238856 239826 238912
rect 240690 228248 240746 228304
rect 240598 164600 240654 164656
rect 240506 153992 240562 154048
rect 240414 138080 240470 138136
rect 241518 85040 241574 85096
rect 241518 74468 241520 74488
rect 241520 74468 241572 74488
rect 241572 74468 241574 74488
rect 241518 74432 241574 74468
rect 241518 58520 241574 58576
rect 242806 233552 242862 233608
rect 242806 222944 242862 223000
rect 242806 217640 242862 217696
rect 241978 212372 241980 212392
rect 241980 212372 242032 212392
rect 242032 212372 242034 212392
rect 241978 212336 242034 212372
rect 242530 207032 242586 207088
rect 242438 201728 242494 201784
rect 242346 196424 242402 196480
rect 241886 191120 241942 191176
rect 242806 185816 242862 185872
rect 242806 180512 242862 180568
rect 242806 175228 242862 175264
rect 242806 175208 242808 175228
rect 242808 175208 242860 175228
rect 242860 175208 242862 175228
rect 241886 169940 241888 169960
rect 241888 169940 241940 169960
rect 241940 169940 241942 169960
rect 241886 169904 241942 169940
rect 241886 159296 241942 159352
rect 242806 148688 242862 148744
rect 241886 143420 241888 143440
rect 241888 143420 241940 143440
rect 241940 143420 241942 143440
rect 241886 143384 241942 143420
rect 242254 127472 242310 127528
rect 241978 122168 242034 122224
rect 242806 116864 242862 116920
rect 241886 111596 241888 111616
rect 241888 111596 241940 111616
rect 241940 111596 241942 111616
rect 241886 111560 241942 111596
rect 241886 106256 241942 106312
rect 241794 100952 241850 101008
rect 242806 95648 242862 95704
rect 242806 90344 242862 90400
rect 242254 79736 242310 79792
rect 241702 69128 241758 69184
rect 242806 63824 242862 63880
rect 241978 53216 242034 53272
rect 241610 47912 241666 47968
rect 240322 42608 240378 42664
rect 243082 132776 243138 132832
rect 337658 376896 337714 376952
rect 337750 375944 337806 376000
rect 337658 373768 337714 373824
rect 337474 372816 337530 372872
rect 337474 371048 337530 371104
rect 337750 369980 337806 370016
rect 337750 369960 337752 369980
rect 337752 369960 337804 369980
rect 337804 369960 337806 369980
rect 337474 368192 337530 368248
rect 337290 349968 337346 350024
rect 337382 348336 337438 348392
rect 337566 348064 337622 348120
rect 267002 244296 267058 244352
rect 356058 338000 356114 338056
rect 368478 338020 368534 338056
rect 368478 338000 368480 338020
rect 368480 338000 368532 338020
rect 368532 338000 368534 338020
rect 371238 338000 371294 338056
rect 382278 338000 382334 338056
rect 386602 338000 386658 338056
rect 407118 338000 407174 338056
rect 363050 337728 363106 337784
rect 367098 337728 367154 337784
rect 356150 337592 356206 337648
rect 357438 337592 357494 337648
rect 358818 337592 358874 337648
rect 360198 337592 360254 337648
rect 362958 337592 363014 337648
rect 361578 337048 361634 337104
rect 364338 337592 364394 337648
rect 365718 337592 365774 337648
rect 367190 337592 367246 337648
rect 378138 337864 378194 337920
rect 371882 337728 371938 337784
rect 376850 337728 376906 337784
rect 371330 337592 371386 337648
rect 369858 336912 369914 336968
rect 369950 336776 370006 336832
rect 370502 38528 370558 38584
rect 372710 337592 372766 337648
rect 373998 337592 374054 337648
rect 376758 337592 376814 337648
rect 375378 337184 375434 337240
rect 375470 337048 375526 337104
rect 379610 337728 379666 337784
rect 379518 337592 379574 337648
rect 380990 337592 381046 337648
rect 380898 337320 380954 337376
rect 383658 337592 383714 337648
rect 385038 337592 385094 337648
rect 382278 337184 382334 337240
rect 385130 337048 385186 337104
rect 386418 337592 386474 337648
rect 391938 337864 391994 337920
rect 394698 337864 394754 337920
rect 396078 337864 396134 337920
rect 398838 337864 398894 337920
rect 387798 337728 387854 337784
rect 390558 337728 390614 337784
rect 387890 337592 387946 337648
rect 389178 337612 389234 337648
rect 389178 337592 389180 337612
rect 389180 337592 389232 337612
rect 389232 337592 389234 337612
rect 390558 337456 390614 337512
rect 393410 337592 393466 337648
rect 392582 336912 392638 336968
rect 393870 337456 393926 337512
rect 396170 337592 396226 337648
rect 397550 337592 397606 337648
rect 397458 337340 397514 337376
rect 397458 337320 397460 337340
rect 397460 337320 397512 337340
rect 397512 337320 397514 337340
rect 402978 337592 403034 337648
rect 405738 337592 405794 337648
rect 400218 336776 400274 336832
rect 409878 337592 409934 337648
rect 412638 337592 412694 337648
rect 415398 337592 415454 337648
rect 417422 337592 417478 337648
rect 420918 337592 420974 337648
rect 424322 337592 424378 337648
rect 427818 337592 427874 337648
rect 430578 337592 430634 337648
rect 433338 337592 433394 337648
rect 440238 337592 440294 337648
rect 442998 337592 443054 337648
rect 422666 336796 422722 336832
rect 422666 336776 422668 336796
rect 422668 336776 422720 336796
rect 422720 336776 422722 336796
rect 434718 337048 434774 337104
rect 437478 337048 437534 337104
rect 445758 337204 445814 337240
rect 445758 337184 445760 337204
rect 445760 337184 445812 337204
rect 445812 337184 445814 337204
rect 580170 697176 580226 697232
rect 580170 683848 580226 683904
rect 580170 670692 580172 670712
rect 580172 670692 580224 670712
rect 580224 670692 580226 670712
rect 580170 670656 580226 670692
rect 580170 644000 580226 644056
rect 580262 630808 580318 630864
rect 580170 617480 580226 617536
rect 580170 590960 580226 591016
rect 580170 577632 580226 577688
rect 580170 564304 580226 564360
rect 579894 537784 579950 537840
rect 580170 524476 580226 524512
rect 580170 524456 580172 524476
rect 580172 524456 580224 524476
rect 580224 524456 580226 524476
rect 580170 511264 580226 511320
rect 580170 484608 580226 484664
rect 580170 458088 580226 458144
rect 580170 418240 580226 418296
rect 580170 404912 580226 404968
rect 580170 365064 580226 365120
rect 580170 351908 580172 351928
rect 580172 351908 580224 351928
rect 580224 351908 580226 351928
rect 580170 351872 580226 351908
rect 580354 471416 580410 471472
rect 580446 431568 580502 431624
rect 580538 378392 580594 378448
rect 580170 325216 580226 325272
rect 580170 312024 580226 312080
rect 580170 298696 580226 298752
rect 579802 272176 579858 272232
rect 580170 258848 580226 258904
rect 579802 245520 579858 245576
rect 579802 232328 579858 232384
rect 579894 205672 579950 205728
rect 580170 192480 580226 192536
rect 580170 165824 580226 165880
rect 579802 152632 579858 152688
rect 580170 139340 580172 139360
rect 580172 139340 580224 139360
rect 580224 139340 580226 139360
rect 580170 139304 580226 139340
rect 580170 125976 580226 126032
rect 580170 112784 580226 112840
rect 580170 99456 580226 99512
rect 580170 86128 580226 86184
rect 579986 72936 580042 72992
rect 580446 219000 580502 219056
rect 580354 179152 580410 179208
rect 580262 59608 580318 59664
rect 580170 46280 580226 46336
rect 580170 33108 580226 33144
rect 580170 33088 580172 33108
rect 580172 33088 580224 33108
rect 580224 33088 580226 33108
rect 580170 19760 580226 19816
rect 580262 6568 580318 6624
<< metal3 >>
rect -960 697220 480 697460
rect 580165 697234 580231 697237
rect 583520 697234 584960 697324
rect 580165 697232 584960 697234
rect 580165 697176 580170 697232
rect 580226 697176 584960 697232
rect 580165 697174 584960 697176
rect 580165 697171 580231 697174
rect 583520 697084 584960 697174
rect -960 684314 480 684404
rect 2773 684314 2839 684317
rect -960 684312 2839 684314
rect -960 684256 2778 684312
rect 2834 684256 2839 684312
rect -960 684254 2839 684256
rect -960 684164 480 684254
rect 2773 684251 2839 684254
rect 580165 683906 580231 683909
rect 583520 683906 584960 683996
rect 580165 683904 584960 683906
rect 580165 683848 580170 683904
rect 580226 683848 584960 683904
rect 580165 683846 584960 683848
rect 580165 683843 580231 683846
rect 583520 683756 584960 683846
rect -960 671258 480 671348
rect 3417 671258 3483 671261
rect -960 671256 3483 671258
rect -960 671200 3422 671256
rect 3478 671200 3483 671256
rect -960 671198 3483 671200
rect -960 671108 480 671198
rect 3417 671195 3483 671198
rect 580165 670714 580231 670717
rect 583520 670714 584960 670804
rect 580165 670712 584960 670714
rect 580165 670656 580170 670712
rect 580226 670656 584960 670712
rect 580165 670654 584960 670656
rect 580165 670651 580231 670654
rect 583520 670564 584960 670654
rect -960 658202 480 658292
rect 3509 658202 3575 658205
rect -960 658200 3575 658202
rect -960 658144 3514 658200
rect 3570 658144 3575 658200
rect -960 658142 3575 658144
rect -960 658052 480 658142
rect 3509 658139 3575 658142
rect 583520 657236 584960 657476
rect -960 644996 480 645236
rect 580165 644058 580231 644061
rect 583520 644058 584960 644148
rect 580165 644056 584960 644058
rect 580165 644000 580170 644056
rect 580226 644000 584960 644056
rect 580165 643998 584960 644000
rect 580165 643995 580231 643998
rect 583520 643908 584960 643998
rect -960 632090 480 632180
rect 3509 632090 3575 632093
rect -960 632088 3575 632090
rect -960 632032 3514 632088
rect 3570 632032 3575 632088
rect -960 632030 3575 632032
rect -960 631940 480 632030
rect 3509 632027 3575 632030
rect 580257 630866 580323 630869
rect 583520 630866 584960 630956
rect 580257 630864 584960 630866
rect 580257 630808 580262 630864
rect 580318 630808 584960 630864
rect 580257 630806 584960 630808
rect 580257 630803 580323 630806
rect 583520 630716 584960 630806
rect -960 619170 480 619260
rect 3509 619170 3575 619173
rect -960 619168 3575 619170
rect -960 619112 3514 619168
rect 3570 619112 3575 619168
rect -960 619110 3575 619112
rect -960 619020 480 619110
rect 3509 619107 3575 619110
rect 580165 617538 580231 617541
rect 583520 617538 584960 617628
rect 580165 617536 584960 617538
rect 580165 617480 580170 617536
rect 580226 617480 584960 617536
rect 580165 617478 584960 617480
rect 580165 617475 580231 617478
rect 583520 617388 584960 617478
rect -960 606114 480 606204
rect 3325 606114 3391 606117
rect -960 606112 3391 606114
rect -960 606056 3330 606112
rect 3386 606056 3391 606112
rect -960 606054 3391 606056
rect -960 605964 480 606054
rect 3325 606051 3391 606054
rect 583520 604060 584960 604300
rect -960 592908 480 593148
rect 580165 591018 580231 591021
rect 583520 591018 584960 591108
rect 580165 591016 584960 591018
rect 580165 590960 580170 591016
rect 580226 590960 584960 591016
rect 580165 590958 584960 590960
rect 580165 590955 580231 590958
rect 583520 590868 584960 590958
rect -960 580002 480 580092
rect 3325 580002 3391 580005
rect -960 580000 3391 580002
rect -960 579944 3330 580000
rect 3386 579944 3391 580000
rect -960 579942 3391 579944
rect -960 579852 480 579942
rect 3325 579939 3391 579942
rect 580165 577690 580231 577693
rect 583520 577690 584960 577780
rect 580165 577688 584960 577690
rect 580165 577632 580170 577688
rect 580226 577632 584960 577688
rect 580165 577630 584960 577632
rect 580165 577627 580231 577630
rect 583520 577540 584960 577630
rect -960 566946 480 567036
rect 3601 566946 3667 566949
rect -960 566944 3667 566946
rect -960 566888 3606 566944
rect 3662 566888 3667 566944
rect -960 566886 3667 566888
rect -960 566796 480 566886
rect 3601 566883 3667 566886
rect 580165 564362 580231 564365
rect 583520 564362 584960 564452
rect 580165 564360 584960 564362
rect 580165 564304 580170 564360
rect 580226 564304 584960 564360
rect 580165 564302 584960 564304
rect 580165 564299 580231 564302
rect 583520 564212 584960 564302
rect -960 553890 480 553980
rect 3325 553890 3391 553893
rect -960 553888 3391 553890
rect -960 553832 3330 553888
rect 3386 553832 3391 553888
rect -960 553830 3391 553832
rect -960 553740 480 553830
rect 3325 553827 3391 553830
rect 583520 551020 584960 551260
rect -960 540684 480 540924
rect 579889 537842 579955 537845
rect 583520 537842 584960 537932
rect 579889 537840 584960 537842
rect 579889 537784 579894 537840
rect 579950 537784 584960 537840
rect 579889 537782 584960 537784
rect 579889 537779 579955 537782
rect 583520 537692 584960 537782
rect -960 527914 480 528004
rect 3325 527914 3391 527917
rect -960 527912 3391 527914
rect -960 527856 3330 527912
rect 3386 527856 3391 527912
rect -960 527854 3391 527856
rect -960 527764 480 527854
rect 3325 527851 3391 527854
rect 580165 524514 580231 524517
rect 583520 524514 584960 524604
rect 580165 524512 584960 524514
rect 580165 524456 580170 524512
rect 580226 524456 584960 524512
rect 580165 524454 584960 524456
rect 580165 524451 580231 524454
rect 583520 524364 584960 524454
rect -960 514858 480 514948
rect 3325 514858 3391 514861
rect -960 514856 3391 514858
rect -960 514800 3330 514856
rect 3386 514800 3391 514856
rect -960 514798 3391 514800
rect -960 514708 480 514798
rect 3325 514795 3391 514798
rect 580165 511322 580231 511325
rect 583520 511322 584960 511412
rect 580165 511320 584960 511322
rect 580165 511264 580170 511320
rect 580226 511264 584960 511320
rect 580165 511262 584960 511264
rect 580165 511259 580231 511262
rect 583520 511172 584960 511262
rect -960 501802 480 501892
rect 2865 501802 2931 501805
rect -960 501800 2931 501802
rect -960 501744 2870 501800
rect 2926 501744 2931 501800
rect -960 501742 2931 501744
rect -960 501652 480 501742
rect 2865 501739 2931 501742
rect 583520 497844 584960 498084
rect -960 488596 480 488836
rect 580165 484666 580231 484669
rect 583520 484666 584960 484756
rect 580165 484664 584960 484666
rect 580165 484608 580170 484664
rect 580226 484608 584960 484664
rect 580165 484606 584960 484608
rect 580165 484603 580231 484606
rect 583520 484516 584960 484606
rect -960 475690 480 475780
rect 3325 475690 3391 475693
rect -960 475688 3391 475690
rect -960 475632 3330 475688
rect 3386 475632 3391 475688
rect -960 475630 3391 475632
rect -960 475540 480 475630
rect 3325 475627 3391 475630
rect 580349 471474 580415 471477
rect 583520 471474 584960 471564
rect 580349 471472 584960 471474
rect 580349 471416 580354 471472
rect 580410 471416 584960 471472
rect 580349 471414 584960 471416
rect 580349 471411 580415 471414
rect 583520 471324 584960 471414
rect -960 462634 480 462724
rect 3325 462634 3391 462637
rect -960 462632 3391 462634
rect -960 462576 3330 462632
rect 3386 462576 3391 462632
rect -960 462574 3391 462576
rect -960 462484 480 462574
rect 3325 462571 3391 462574
rect 580165 458146 580231 458149
rect 583520 458146 584960 458236
rect 580165 458144 584960 458146
rect 580165 458088 580170 458144
rect 580226 458088 584960 458144
rect 580165 458086 584960 458088
rect 580165 458083 580231 458086
rect 583520 457996 584960 458086
rect -960 449578 480 449668
rect 3325 449578 3391 449581
rect -960 449576 3391 449578
rect -960 449520 3330 449576
rect 3386 449520 3391 449576
rect -960 449518 3391 449520
rect -960 449428 480 449518
rect 3325 449515 3391 449518
rect 583520 444668 584960 444908
rect -960 436508 480 436748
rect 580441 431626 580507 431629
rect 583520 431626 584960 431716
rect 580441 431624 584960 431626
rect 580441 431568 580446 431624
rect 580502 431568 584960 431624
rect 580441 431566 584960 431568
rect 580441 431563 580507 431566
rect 583520 431476 584960 431566
rect -960 423602 480 423692
rect 3141 423602 3207 423605
rect -960 423600 3207 423602
rect -960 423544 3146 423600
rect 3202 423544 3207 423600
rect -960 423542 3207 423544
rect -960 423452 480 423542
rect 3141 423539 3207 423542
rect 580165 418298 580231 418301
rect 583520 418298 584960 418388
rect 580165 418296 584960 418298
rect 580165 418240 580170 418296
rect 580226 418240 584960 418296
rect 580165 418238 584960 418240
rect 580165 418235 580231 418238
rect 583520 418148 584960 418238
rect -960 410546 480 410636
rect 3693 410546 3759 410549
rect -960 410544 3759 410546
rect -960 410488 3698 410544
rect 3754 410488 3759 410544
rect -960 410486 3759 410488
rect -960 410396 480 410486
rect 3693 410483 3759 410486
rect 580165 404970 580231 404973
rect 583520 404970 584960 405060
rect 580165 404968 584960 404970
rect 580165 404912 580170 404968
rect 580226 404912 584960 404968
rect 580165 404910 584960 404912
rect 580165 404907 580231 404910
rect 583520 404820 584960 404910
rect -960 397490 480 397580
rect 3325 397490 3391 397493
rect -960 397488 3391 397490
rect -960 397432 3330 397488
rect 3386 397432 3391 397488
rect -960 397430 3391 397432
rect -960 397340 480 397430
rect 3325 397427 3391 397430
rect 583520 391628 584960 391868
rect -960 384284 480 384524
rect 580533 378450 580599 378453
rect 583520 378450 584960 378540
rect 580533 378448 584960 378450
rect 580533 378392 580538 378448
rect 580594 378392 584960 378448
rect 580533 378390 584960 378392
rect 580533 378387 580599 378390
rect 583520 378300 584960 378390
rect 38469 376954 38535 376957
rect 337653 376954 337719 376957
rect 38469 376952 39498 376954
rect 38469 376896 38474 376952
rect 38530 376924 39498 376952
rect 337653 376952 339418 376954
rect 38530 376896 40020 376924
rect 38469 376894 40020 376896
rect 38469 376891 38535 376894
rect 39438 376864 40020 376894
rect 337653 376896 337658 376952
rect 337714 376924 339418 376952
rect 337714 376896 340032 376924
rect 337653 376894 340032 376896
rect 337653 376891 337719 376894
rect 339358 376864 340032 376894
rect 37917 376002 37983 376005
rect 337745 376002 337811 376005
rect 37917 376000 39498 376002
rect 37917 375944 37922 376000
rect 37978 375972 39498 376000
rect 337745 376000 339418 376002
rect 37978 375944 40020 375972
rect 37917 375942 40020 375944
rect 37917 375939 37983 375942
rect 39438 375912 40020 375942
rect 337745 375944 337750 376000
rect 337806 375972 339418 376000
rect 337806 375944 340032 375972
rect 337745 375942 340032 375944
rect 337745 375939 337811 375942
rect 339358 375912 340032 375942
rect 38101 373826 38167 373829
rect 337653 373826 337719 373829
rect 38101 373824 39498 373826
rect 38101 373768 38106 373824
rect 38162 373796 39498 373824
rect 337653 373824 339418 373826
rect 38162 373768 40020 373796
rect 38101 373766 40020 373768
rect 38101 373763 38167 373766
rect 39438 373736 40020 373766
rect 337653 373768 337658 373824
rect 337714 373796 339418 373824
rect 337714 373768 340032 373796
rect 337653 373766 340032 373768
rect 337653 373763 337719 373766
rect 339358 373736 340032 373766
rect 38285 372874 38351 372877
rect 337469 372874 337535 372877
rect 38285 372872 39498 372874
rect 38285 372816 38290 372872
rect 38346 372844 39498 372872
rect 337469 372872 339418 372874
rect 38346 372816 40020 372844
rect 38285 372814 40020 372816
rect 38285 372811 38351 372814
rect 39438 372784 40020 372814
rect 337469 372816 337474 372872
rect 337530 372844 339418 372872
rect 337530 372816 340032 372844
rect 337469 372814 340032 372816
rect 337469 372811 337535 372814
rect 339358 372784 340032 372814
rect -960 371378 480 371468
rect 3325 371378 3391 371381
rect -960 371376 3391 371378
rect -960 371320 3330 371376
rect 3386 371320 3391 371376
rect -960 371318 3391 371320
rect -960 371228 480 371318
rect 3325 371315 3391 371318
rect 38837 371106 38903 371109
rect 337469 371106 337535 371109
rect 38837 371104 39498 371106
rect 38837 371048 38842 371104
rect 38898 371076 39498 371104
rect 337469 371104 339418 371106
rect 38898 371048 40020 371076
rect 38837 371046 40020 371048
rect 38837 371043 38903 371046
rect 39438 371016 40020 371046
rect 337469 371048 337474 371104
rect 337530 371076 339418 371104
rect 337530 371048 340032 371076
rect 337469 371046 340032 371048
rect 337469 371043 337535 371046
rect 339358 371016 340032 371046
rect 38653 370018 38719 370021
rect 337745 370018 337811 370021
rect 38653 370016 39498 370018
rect 38653 369960 38658 370016
rect 38714 369988 39498 370016
rect 337745 370016 339418 370018
rect 38714 369960 40020 369988
rect 38653 369958 40020 369960
rect 38653 369955 38719 369958
rect 39438 369928 40020 369958
rect 337745 369960 337750 370016
rect 337806 369988 339418 370016
rect 337806 369960 340032 369988
rect 337745 369958 340032 369960
rect 337745 369955 337811 369958
rect 339358 369928 340032 369958
rect 38745 368250 38811 368253
rect 337469 368250 337535 368253
rect 38745 368248 39498 368250
rect 38745 368192 38750 368248
rect 38806 368220 39498 368248
rect 337469 368248 339418 368250
rect 38806 368192 40020 368220
rect 38745 368190 40020 368192
rect 38745 368187 38811 368190
rect 39438 368160 40020 368190
rect 337469 368192 337474 368248
rect 337530 368220 339418 368248
rect 337530 368192 340032 368220
rect 337469 368190 340032 368192
rect 337469 368187 337535 368190
rect 339358 368160 340032 368190
rect 580165 365122 580231 365125
rect 583520 365122 584960 365212
rect 580165 365120 584960 365122
rect 580165 365064 580170 365120
rect 580226 365064 584960 365120
rect 580165 365062 584960 365064
rect 580165 365059 580231 365062
rect 583520 364972 584960 365062
rect -960 358458 480 358548
rect 3785 358458 3851 358461
rect -960 358456 3851 358458
rect -960 358400 3790 358456
rect 3846 358400 3851 358456
rect -960 358398 3851 358400
rect -960 358308 480 358398
rect 3785 358395 3851 358398
rect 580165 351930 580231 351933
rect 583520 351930 584960 352020
rect 580165 351928 584960 351930
rect 580165 351872 580170 351928
rect 580226 351872 584960 351928
rect 580165 351870 584960 351872
rect 580165 351867 580231 351870
rect 583520 351780 584960 351870
rect 38377 350026 38443 350029
rect 337285 350026 337351 350029
rect 38377 350024 39498 350026
rect 38377 349968 38382 350024
rect 38438 349996 39498 350024
rect 337285 350024 339418 350026
rect 38438 349968 40020 349996
rect 38377 349966 40020 349968
rect 38377 349963 38443 349966
rect 39438 349936 40020 349966
rect 337285 349968 337290 350024
rect 337346 349996 339418 350024
rect 337346 349968 340032 349996
rect 337285 349966 340032 349968
rect 337285 349963 337351 349966
rect 339358 349936 340032 349966
rect 38561 348394 38627 348397
rect 337377 348394 337443 348397
rect 38561 348392 39498 348394
rect 38561 348336 38566 348392
rect 38622 348364 39498 348392
rect 337377 348392 339418 348394
rect 38622 348336 40020 348364
rect 38561 348334 40020 348336
rect 38561 348331 38627 348334
rect 39438 348304 40020 348334
rect 337377 348336 337382 348392
rect 337438 348364 339418 348392
rect 337438 348336 340032 348364
rect 337377 348334 340032 348336
rect 337377 348331 337443 348334
rect 339358 348304 340032 348334
rect 37825 348122 37891 348125
rect 337561 348122 337627 348125
rect 37825 348120 39498 348122
rect 37825 348064 37830 348120
rect 37886 348092 39498 348120
rect 337561 348120 339418 348122
rect 37886 348064 40020 348092
rect 37825 348062 40020 348064
rect 37825 348059 37891 348062
rect 39438 348032 40020 348062
rect 337561 348064 337566 348120
rect 337622 348092 339418 348120
rect 337622 348064 340032 348092
rect 337561 348062 340032 348064
rect 337561 348059 337627 348062
rect 339358 348032 340032 348062
rect -960 345402 480 345492
rect 3049 345402 3115 345405
rect -960 345400 3115 345402
rect -960 345344 3054 345400
rect 3110 345344 3115 345400
rect -960 345342 3115 345344
rect -960 345252 480 345342
rect 3049 345339 3115 345342
rect 583520 338452 584960 338692
rect 76966 338132 76972 338196
rect 77036 338132 77042 338196
rect 90950 338132 90956 338196
rect 91020 338132 91026 338196
rect 131062 338132 131068 338196
rect 131132 338132 131138 338196
rect 372286 338132 372292 338196
rect 372356 338132 372362 338196
rect 382774 338132 382780 338196
rect 382844 338132 382850 338196
rect 386454 338132 386460 338196
rect 386524 338132 386530 338196
rect 408166 338132 408172 338196
rect 408236 338132 408242 338196
rect 76281 338058 76347 338061
rect 76974 338058 77034 338132
rect 76281 338056 77034 338058
rect 76281 338000 76286 338056
rect 76342 338000 77034 338056
rect 76281 337998 77034 338000
rect 90958 338061 91018 338132
rect 131070 338061 131130 338132
rect 90958 338056 91067 338061
rect 90958 338000 91006 338056
rect 91062 338000 91067 338056
rect 90958 337998 91067 338000
rect 76281 337995 76347 337998
rect 91001 337995 91067 337998
rect 131021 338056 131130 338061
rect 356053 338060 356119 338061
rect 356053 338058 356100 338060
rect 131021 338000 131026 338056
rect 131082 338000 131130 338056
rect 131021 337998 131130 338000
rect 356008 338056 356100 338058
rect 356008 338000 356058 338056
rect 356008 337998 356100 338000
rect 131021 337995 131087 337998
rect 356053 337996 356100 337998
rect 356164 337996 356170 338060
rect 368473 338058 368539 338061
rect 368974 338058 368980 338060
rect 368473 338056 368980 338058
rect 368473 338000 368478 338056
rect 368534 338000 368980 338056
rect 368473 337998 368980 338000
rect 356053 337995 356119 337996
rect 368473 337995 368539 337998
rect 368974 337996 368980 337998
rect 369044 337996 369050 338060
rect 371233 338058 371299 338061
rect 372294 338058 372354 338132
rect 371233 338056 372354 338058
rect 371233 338000 371238 338056
rect 371294 338000 372354 338056
rect 371233 337998 372354 338000
rect 382273 338058 382339 338061
rect 382782 338058 382842 338132
rect 382273 338056 382842 338058
rect 382273 338000 382278 338056
rect 382334 338000 382842 338056
rect 382273 337998 382842 338000
rect 386462 338058 386522 338132
rect 386597 338058 386663 338061
rect 386462 338056 386663 338058
rect 386462 338000 386602 338056
rect 386658 338000 386663 338056
rect 386462 337998 386663 338000
rect 371233 337995 371299 337998
rect 382273 337995 382339 337998
rect 386597 337995 386663 337998
rect 407113 338058 407179 338061
rect 408174 338058 408234 338132
rect 407113 338056 408234 338058
rect 407113 338000 407118 338056
rect 407174 338000 408234 338056
rect 407113 337998 408234 338000
rect 407113 337995 407179 337998
rect 55990 337860 55996 337924
rect 56060 337922 56066 337924
rect 56501 337922 56567 337925
rect 68318 337922 68324 337924
rect 56060 337920 56567 337922
rect 56060 337864 56506 337920
rect 56562 337864 56567 337920
rect 56060 337862 56567 337864
rect 56060 337860 56066 337862
rect 56501 337859 56567 337862
rect 64830 337862 68324 337922
rect 47710 337724 47716 337788
rect 47780 337786 47786 337788
rect 64830 337786 64890 337862
rect 68318 337860 68324 337862
rect 68388 337860 68394 337924
rect 78070 337860 78076 337924
rect 78140 337922 78146 337924
rect 78581 337922 78647 337925
rect 78140 337920 78647 337922
rect 78140 337864 78586 337920
rect 78642 337864 78647 337920
rect 78140 337862 78647 337864
rect 78140 337860 78146 337862
rect 78581 337859 78647 337862
rect 97942 337860 97948 337924
rect 98012 337922 98018 337924
rect 99281 337922 99347 337925
rect 98012 337920 99347 337922
rect 98012 337864 99286 337920
rect 99342 337864 99347 337920
rect 98012 337862 99347 337864
rect 98012 337860 98018 337862
rect 99281 337859 99347 337862
rect 378133 337922 378199 337925
rect 378542 337922 378548 337924
rect 378133 337920 378548 337922
rect 378133 337864 378138 337920
rect 378194 337864 378548 337920
rect 378133 337862 378548 337864
rect 378133 337859 378199 337862
rect 378542 337860 378548 337862
rect 378612 337860 378618 337924
rect 391933 337922 391999 337925
rect 392158 337922 392164 337924
rect 391933 337920 392164 337922
rect 391933 337864 391938 337920
rect 391994 337864 392164 337920
rect 391933 337862 392164 337864
rect 391933 337859 391999 337862
rect 392158 337860 392164 337862
rect 392228 337860 392234 337924
rect 394693 337922 394759 337925
rect 395654 337922 395660 337924
rect 394693 337920 395660 337922
rect 394693 337864 394698 337920
rect 394754 337864 395660 337920
rect 394693 337862 395660 337864
rect 394693 337859 394759 337862
rect 395654 337860 395660 337862
rect 395724 337860 395730 337924
rect 396073 337922 396139 337925
rect 396574 337922 396580 337924
rect 396073 337920 396580 337922
rect 396073 337864 396078 337920
rect 396134 337864 396580 337920
rect 396073 337862 396580 337864
rect 396073 337859 396139 337862
rect 396574 337860 396580 337862
rect 396644 337860 396650 337924
rect 398833 337922 398899 337925
rect 399150 337922 399156 337924
rect 398833 337920 399156 337922
rect 398833 337864 398838 337920
rect 398894 337864 399156 337920
rect 398833 337862 399156 337864
rect 398833 337859 398899 337862
rect 399150 337860 399156 337862
rect 399220 337860 399226 337924
rect 47780 337726 64890 337786
rect 47780 337724 47786 337726
rect 67582 337724 67588 337788
rect 67652 337786 67658 337788
rect 68921 337786 68987 337789
rect 67652 337784 68987 337786
rect 67652 337728 68926 337784
rect 68982 337728 68987 337784
rect 67652 337726 68987 337728
rect 67652 337724 67658 337726
rect 68921 337723 68987 337726
rect 70577 337786 70643 337789
rect 71262 337786 71268 337788
rect 70577 337784 71268 337786
rect 70577 337728 70582 337784
rect 70638 337728 71268 337784
rect 70577 337726 71268 337728
rect 70577 337723 70643 337726
rect 71262 337724 71268 337726
rect 71332 337724 71338 337788
rect 73470 337724 73476 337788
rect 73540 337786 73546 337788
rect 74349 337786 74415 337789
rect 73540 337784 74415 337786
rect 73540 337728 74354 337784
rect 74410 337728 74415 337784
rect 73540 337726 74415 337728
rect 73540 337724 73546 337726
rect 74349 337723 74415 337726
rect 75862 337724 75868 337788
rect 75932 337786 75938 337788
rect 77201 337786 77267 337789
rect 75932 337784 77267 337786
rect 75932 337728 77206 337784
rect 77262 337728 77267 337784
rect 75932 337726 77267 337728
rect 75932 337724 75938 337726
rect 77201 337723 77267 337726
rect 82854 337724 82860 337788
rect 82924 337786 82930 337788
rect 83549 337786 83615 337789
rect 82924 337784 83615 337786
rect 82924 337728 83554 337784
rect 83610 337728 83615 337784
rect 82924 337726 83615 337728
rect 82924 337724 82930 337726
rect 83549 337723 83615 337726
rect 87638 337724 87644 337788
rect 87708 337786 87714 337788
rect 88057 337786 88123 337789
rect 87708 337784 88123 337786
rect 87708 337728 88062 337784
rect 88118 337728 88123 337784
rect 87708 337726 88123 337728
rect 87708 337724 87714 337726
rect 88057 337723 88123 337726
rect 91502 337724 91508 337788
rect 91572 337786 91578 337788
rect 92381 337786 92447 337789
rect 91572 337784 92447 337786
rect 91572 337728 92386 337784
rect 92442 337728 92447 337784
rect 91572 337726 92447 337728
rect 91572 337724 91578 337726
rect 92381 337723 92447 337726
rect 93342 337724 93348 337788
rect 93412 337786 93418 337788
rect 93577 337786 93643 337789
rect 93412 337784 93643 337786
rect 93412 337728 93582 337784
rect 93638 337728 93643 337784
rect 93412 337726 93643 337728
rect 93412 337724 93418 337726
rect 93577 337723 93643 337726
rect 94262 337724 94268 337788
rect 94332 337786 94338 337788
rect 95141 337786 95207 337789
rect 94332 337784 95207 337786
rect 94332 337728 95146 337784
rect 95202 337728 95207 337784
rect 94332 337726 95207 337728
rect 94332 337724 94338 337726
rect 95141 337723 95207 337726
rect 97993 337786 98059 337789
rect 99046 337786 99052 337788
rect 97993 337784 99052 337786
rect 97993 337728 97998 337784
rect 98054 337728 99052 337784
rect 97993 337726 99052 337728
rect 97993 337723 98059 337726
rect 99046 337724 99052 337726
rect 99116 337724 99122 337788
rect 142153 337786 142219 337789
rect 143390 337786 143396 337788
rect 142153 337784 143396 337786
rect 142153 337728 142158 337784
rect 142214 337728 143396 337784
rect 142153 337726 143396 337728
rect 142153 337723 142219 337726
rect 143390 337724 143396 337726
rect 143460 337724 143466 337788
rect 363045 337786 363111 337789
rect 364190 337786 364196 337788
rect 363045 337784 364196 337786
rect 363045 337728 363050 337784
rect 363106 337728 364196 337784
rect 363045 337726 364196 337728
rect 363045 337723 363111 337726
rect 364190 337724 364196 337726
rect 364260 337724 364266 337788
rect 367093 337786 367159 337789
rect 368054 337786 368060 337788
rect 367093 337784 368060 337786
rect 367093 337728 367098 337784
rect 367154 337728 368060 337784
rect 367093 337726 368060 337728
rect 367093 337723 367159 337726
rect 368054 337724 368060 337726
rect 368124 337724 368130 337788
rect 371877 337786 371943 337789
rect 373574 337786 373580 337788
rect 371877 337784 373580 337786
rect 371877 337728 371882 337784
rect 371938 337728 373580 337784
rect 371877 337726 373580 337728
rect 371877 337723 371943 337726
rect 373574 337724 373580 337726
rect 373644 337724 373650 337788
rect 376845 337786 376911 337789
rect 377990 337786 377996 337788
rect 376845 337784 377996 337786
rect 376845 337728 376850 337784
rect 376906 337728 377996 337784
rect 376845 337726 377996 337728
rect 376845 337723 376911 337726
rect 377990 337724 377996 337726
rect 378060 337724 378066 337788
rect 379605 337786 379671 337789
rect 380566 337786 380572 337788
rect 379605 337784 380572 337786
rect 379605 337728 379610 337784
rect 379666 337728 380572 337784
rect 379605 337726 380572 337728
rect 379605 337723 379671 337726
rect 380566 337724 380572 337726
rect 380636 337724 380642 337788
rect 387793 337786 387859 337789
rect 388662 337786 388668 337788
rect 387793 337784 388668 337786
rect 387793 337728 387798 337784
rect 387854 337728 388668 337784
rect 387793 337726 388668 337728
rect 387793 337723 387859 337726
rect 388662 337724 388668 337726
rect 388732 337724 388738 337788
rect 390553 337786 390619 337789
rect 391054 337786 391060 337788
rect 390553 337784 391060 337786
rect 390553 337728 390558 337784
rect 390614 337728 391060 337784
rect 390553 337726 391060 337728
rect 390553 337723 390619 337726
rect 391054 337724 391060 337726
rect 391124 337724 391130 337788
rect 58198 337588 58204 337652
rect 58268 337650 58274 337652
rect 59261 337650 59327 337653
rect 58268 337648 59327 337650
rect 58268 337592 59266 337648
rect 59322 337592 59327 337648
rect 58268 337590 59327 337592
rect 58268 337588 58274 337590
rect 59261 337587 59327 337590
rect 61878 337588 61884 337652
rect 61948 337650 61954 337652
rect 62021 337650 62087 337653
rect 61948 337648 62087 337650
rect 61948 337592 62026 337648
rect 62082 337592 62087 337648
rect 61948 337590 62087 337592
rect 61948 337588 61954 337590
rect 62021 337587 62087 337590
rect 63166 337588 63172 337652
rect 63236 337650 63242 337652
rect 63401 337650 63467 337653
rect 63236 337648 63467 337650
rect 63236 337592 63406 337648
rect 63462 337592 63467 337648
rect 63236 337590 63467 337592
rect 63236 337588 63242 337590
rect 63401 337587 63467 337590
rect 64965 337650 65031 337653
rect 65374 337650 65380 337652
rect 64965 337648 65380 337650
rect 64965 337592 64970 337648
rect 65026 337592 65380 337648
rect 64965 337590 65380 337592
rect 64965 337587 65031 337590
rect 65374 337588 65380 337590
rect 65444 337588 65450 337652
rect 66345 337650 66411 337653
rect 66662 337650 66668 337652
rect 66345 337648 66668 337650
rect 66345 337592 66350 337648
rect 66406 337592 66668 337648
rect 66345 337590 66668 337592
rect 66345 337587 66411 337590
rect 66662 337588 66668 337590
rect 66732 337588 66738 337652
rect 67633 337650 67699 337653
rect 68686 337650 68692 337652
rect 67633 337648 68692 337650
rect 67633 337592 67638 337648
rect 67694 337592 68692 337648
rect 67633 337590 68692 337592
rect 67633 337587 67699 337590
rect 68686 337588 68692 337590
rect 68756 337588 68762 337652
rect 70485 337650 70551 337653
rect 70710 337650 70716 337652
rect 70485 337648 70716 337650
rect 70485 337592 70490 337648
rect 70546 337592 70716 337648
rect 70485 337590 70716 337592
rect 70485 337587 70551 337590
rect 70710 337588 70716 337590
rect 70780 337588 70786 337652
rect 73654 337588 73660 337652
rect 73724 337650 73730 337652
rect 74441 337650 74507 337653
rect 73724 337648 74507 337650
rect 73724 337592 74446 337648
rect 74502 337592 74507 337648
rect 73724 337590 74507 337592
rect 73724 337588 73730 337590
rect 74441 337587 74507 337590
rect 74574 337588 74580 337652
rect 74644 337650 74650 337652
rect 74901 337650 74967 337653
rect 78489 337652 78555 337653
rect 74644 337648 74967 337650
rect 74644 337592 74906 337648
rect 74962 337592 74967 337648
rect 74644 337590 74967 337592
rect 74644 337588 74650 337590
rect 74901 337587 74967 337590
rect 78438 337588 78444 337652
rect 78508 337650 78555 337652
rect 78508 337648 78600 337650
rect 78550 337592 78600 337648
rect 78508 337590 78600 337592
rect 78508 337588 78555 337590
rect 79542 337588 79548 337652
rect 79612 337650 79618 337652
rect 79961 337650 80027 337653
rect 81065 337652 81131 337653
rect 79612 337648 80027 337650
rect 79612 337592 79966 337648
rect 80022 337592 80027 337648
rect 79612 337590 80027 337592
rect 79612 337588 79618 337590
rect 78489 337587 78555 337588
rect 79961 337587 80027 337590
rect 81014 337588 81020 337652
rect 81084 337650 81131 337652
rect 81084 337648 81176 337650
rect 81126 337592 81176 337648
rect 81084 337590 81176 337592
rect 81084 337588 81131 337590
rect 81750 337588 81756 337652
rect 81820 337650 81826 337652
rect 82721 337650 82787 337653
rect 81820 337648 82787 337650
rect 81820 337592 82726 337648
rect 82782 337592 82787 337648
rect 81820 337590 82787 337592
rect 81820 337588 81826 337590
rect 81065 337587 81131 337588
rect 82721 337587 82787 337590
rect 82905 337650 82971 337653
rect 85297 337652 85363 337653
rect 86401 337652 86467 337653
rect 83406 337650 83412 337652
rect 82905 337648 83412 337650
rect 82905 337592 82910 337648
rect 82966 337592 83412 337648
rect 82905 337590 83412 337592
rect 82905 337587 82971 337590
rect 83406 337588 83412 337590
rect 83476 337588 83482 337652
rect 85246 337588 85252 337652
rect 85316 337650 85363 337652
rect 85316 337648 85408 337650
rect 85358 337592 85408 337648
rect 85316 337590 85408 337592
rect 85316 337588 85363 337590
rect 86350 337588 86356 337652
rect 86420 337650 86467 337652
rect 88149 337652 88215 337653
rect 88149 337650 88196 337652
rect 86420 337648 86512 337650
rect 86462 337592 86512 337648
rect 86420 337590 86512 337592
rect 88104 337648 88196 337650
rect 88104 337592 88154 337648
rect 88104 337590 88196 337592
rect 86420 337588 86467 337590
rect 85297 337587 85363 337588
rect 86401 337587 86467 337588
rect 88149 337588 88196 337590
rect 88260 337588 88266 337652
rect 88425 337650 88491 337653
rect 88742 337650 88748 337652
rect 88425 337648 88748 337650
rect 88425 337592 88430 337648
rect 88486 337592 88748 337648
rect 88425 337590 88748 337592
rect 88149 337587 88215 337588
rect 88425 337587 88491 337590
rect 88742 337588 88748 337590
rect 88812 337588 88818 337652
rect 89846 337588 89852 337652
rect 89916 337650 89922 337652
rect 90633 337650 90699 337653
rect 89916 337648 90699 337650
rect 89916 337592 90638 337648
rect 90694 337592 90699 337648
rect 89916 337590 90699 337592
rect 89916 337588 89922 337590
rect 90633 337587 90699 337590
rect 91185 337650 91251 337653
rect 92238 337650 92244 337652
rect 91185 337648 92244 337650
rect 91185 337592 91190 337648
rect 91246 337592 92244 337648
rect 91185 337590 92244 337592
rect 91185 337587 91251 337590
rect 92238 337588 92244 337590
rect 92308 337588 92314 337652
rect 92473 337650 92539 337653
rect 93526 337650 93532 337652
rect 92473 337648 93532 337650
rect 92473 337592 92478 337648
rect 92534 337592 93532 337648
rect 92473 337590 93532 337592
rect 92473 337587 92539 337590
rect 93526 337588 93532 337590
rect 93596 337588 93602 337652
rect 95734 337588 95740 337652
rect 95804 337650 95810 337652
rect 96337 337650 96403 337653
rect 95804 337648 96403 337650
rect 95804 337592 96342 337648
rect 96398 337592 96403 337648
rect 95804 337590 96403 337592
rect 95804 337588 95810 337590
rect 96337 337587 96403 337590
rect 97022 337588 97028 337652
rect 97092 337650 97098 337652
rect 97901 337650 97967 337653
rect 97092 337648 97967 337650
rect 97092 337592 97906 337648
rect 97962 337592 97967 337648
rect 97092 337590 97967 337592
rect 97092 337588 97098 337590
rect 97901 337587 97967 337590
rect 100753 337650 100819 337653
rect 100886 337650 100892 337652
rect 100753 337648 100892 337650
rect 100753 337592 100758 337648
rect 100814 337592 100892 337648
rect 100753 337590 100892 337592
rect 100753 337587 100819 337590
rect 100886 337588 100892 337590
rect 100956 337588 100962 337652
rect 106038 337588 106044 337652
rect 106108 337650 106114 337652
rect 106181 337650 106247 337653
rect 106108 337648 106247 337650
rect 106108 337592 106186 337648
rect 106242 337592 106247 337648
rect 106108 337590 106247 337592
rect 106108 337588 106114 337590
rect 106181 337587 106247 337590
rect 107653 337650 107719 337653
rect 108246 337650 108252 337652
rect 107653 337648 108252 337650
rect 107653 337592 107658 337648
rect 107714 337592 108252 337648
rect 107653 337590 108252 337592
rect 107653 337587 107719 337590
rect 108246 337588 108252 337590
rect 108316 337588 108322 337652
rect 111006 337588 111012 337652
rect 111076 337650 111082 337652
rect 111701 337650 111767 337653
rect 111076 337648 111767 337650
rect 111076 337592 111706 337648
rect 111762 337592 111767 337648
rect 111076 337590 111767 337592
rect 111076 337588 111082 337590
rect 111701 337587 111767 337590
rect 113173 337650 113239 337653
rect 118601 337652 118667 337653
rect 113398 337650 113404 337652
rect 113173 337648 113404 337650
rect 113173 337592 113178 337648
rect 113234 337592 113404 337648
rect 113173 337590 113404 337592
rect 113173 337587 113239 337590
rect 113398 337588 113404 337590
rect 113468 337588 113474 337652
rect 118550 337588 118556 337652
rect 118620 337650 118667 337652
rect 118620 337648 118712 337650
rect 118662 337592 118712 337648
rect 118620 337590 118712 337592
rect 118620 337588 118667 337590
rect 120942 337588 120948 337652
rect 121012 337650 121018 337652
rect 121361 337650 121427 337653
rect 121012 337648 121427 337650
rect 121012 337592 121366 337648
rect 121422 337592 121427 337648
rect 121012 337590 121427 337592
rect 121012 337588 121018 337590
rect 118601 337587 118667 337588
rect 121361 337587 121427 337590
rect 122833 337650 122899 337653
rect 123518 337650 123524 337652
rect 122833 337648 123524 337650
rect 122833 337592 122838 337648
rect 122894 337592 123524 337648
rect 122833 337590 123524 337592
rect 122833 337587 122899 337590
rect 123518 337588 123524 337590
rect 123588 337588 123594 337652
rect 125910 337588 125916 337652
rect 125980 337650 125986 337652
rect 126881 337650 126947 337653
rect 125980 337648 126947 337650
rect 125980 337592 126886 337648
rect 126942 337592 126947 337648
rect 125980 337590 126947 337592
rect 125980 337588 125986 337590
rect 126881 337587 126947 337590
rect 128486 337588 128492 337652
rect 128556 337650 128562 337652
rect 129641 337650 129707 337653
rect 128556 337648 129707 337650
rect 128556 337592 129646 337648
rect 129702 337592 129707 337648
rect 128556 337590 129707 337592
rect 128556 337588 128562 337590
rect 129641 337587 129707 337590
rect 132585 337650 132651 337653
rect 133454 337650 133460 337652
rect 132585 337648 133460 337650
rect 132585 337592 132590 337648
rect 132646 337592 133460 337648
rect 132585 337590 133460 337592
rect 132585 337587 132651 337590
rect 133454 337588 133460 337590
rect 133524 337588 133530 337652
rect 135253 337650 135319 337653
rect 135846 337650 135852 337652
rect 135253 337648 135852 337650
rect 135253 337592 135258 337648
rect 135314 337592 135852 337648
rect 135253 337590 135852 337592
rect 135253 337587 135319 337590
rect 135846 337588 135852 337590
rect 135916 337588 135922 337652
rect 138606 337588 138612 337652
rect 138676 337650 138682 337652
rect 139301 337650 139367 337653
rect 138676 337648 139367 337650
rect 138676 337592 139306 337648
rect 139362 337592 139367 337648
rect 138676 337590 139367 337592
rect 138676 337588 138682 337590
rect 139301 337587 139367 337590
rect 140998 337588 141004 337652
rect 141068 337650 141074 337652
rect 142061 337650 142127 337653
rect 141068 337648 142127 337650
rect 141068 337592 142066 337648
rect 142122 337592 142127 337648
rect 141068 337590 142127 337592
rect 141068 337588 141074 337590
rect 142061 337587 142127 337590
rect 145966 337588 145972 337652
rect 146036 337650 146042 337652
rect 146201 337650 146267 337653
rect 146036 337648 146267 337650
rect 146036 337592 146206 337648
rect 146262 337592 146267 337648
rect 146036 337590 146267 337592
rect 146036 337588 146042 337590
rect 146201 337587 146267 337590
rect 356145 337650 356211 337653
rect 357014 337650 357020 337652
rect 356145 337648 357020 337650
rect 356145 337592 356150 337648
rect 356206 337592 357020 337648
rect 356145 337590 357020 337592
rect 356145 337587 356211 337590
rect 357014 337588 357020 337590
rect 357084 337588 357090 337652
rect 357433 337650 357499 337653
rect 358118 337650 358124 337652
rect 357433 337648 358124 337650
rect 357433 337592 357438 337648
rect 357494 337592 358124 337648
rect 357433 337590 358124 337592
rect 357433 337587 357499 337590
rect 358118 337588 358124 337590
rect 358188 337588 358194 337652
rect 358813 337650 358879 337653
rect 359590 337650 359596 337652
rect 358813 337648 359596 337650
rect 358813 337592 358818 337648
rect 358874 337592 359596 337648
rect 358813 337590 359596 337592
rect 358813 337587 358879 337590
rect 359590 337588 359596 337590
rect 359660 337588 359666 337652
rect 360193 337650 360259 337653
rect 360510 337650 360516 337652
rect 360193 337648 360516 337650
rect 360193 337592 360198 337648
rect 360254 337592 360516 337648
rect 360193 337590 360516 337592
rect 360193 337587 360259 337590
rect 360510 337588 360516 337590
rect 360580 337588 360586 337652
rect 362953 337650 363019 337653
rect 363086 337650 363092 337652
rect 362953 337648 363092 337650
rect 362953 337592 362958 337648
rect 363014 337592 363092 337648
rect 362953 337590 363092 337592
rect 362953 337587 363019 337590
rect 363086 337588 363092 337590
rect 363156 337588 363162 337652
rect 364333 337650 364399 337653
rect 365478 337650 365484 337652
rect 364333 337648 365484 337650
rect 364333 337592 364338 337648
rect 364394 337592 365484 337648
rect 364333 337590 365484 337592
rect 364333 337587 364399 337590
rect 365478 337588 365484 337590
rect 365548 337588 365554 337652
rect 365713 337650 365779 337653
rect 366398 337650 366404 337652
rect 365713 337648 366404 337650
rect 365713 337592 365718 337648
rect 365774 337592 366404 337648
rect 365713 337590 366404 337592
rect 365713 337587 365779 337590
rect 366398 337588 366404 337590
rect 366468 337588 366474 337652
rect 367185 337650 367251 337653
rect 371325 337652 371391 337653
rect 367502 337650 367508 337652
rect 367185 337648 367508 337650
rect 367185 337592 367190 337648
rect 367246 337592 367508 337648
rect 367185 337590 367508 337592
rect 367185 337587 367251 337590
rect 367502 337588 367508 337590
rect 367572 337588 367578 337652
rect 371325 337650 371372 337652
rect 371280 337648 371372 337650
rect 371280 337592 371330 337648
rect 371280 337590 371372 337592
rect 371325 337588 371372 337590
rect 371436 337588 371442 337652
rect 372705 337650 372771 337653
rect 373390 337650 373396 337652
rect 372705 337648 373396 337650
rect 372705 337592 372710 337648
rect 372766 337592 373396 337648
rect 372705 337590 373396 337592
rect 371325 337587 371391 337588
rect 372705 337587 372771 337590
rect 373390 337588 373396 337590
rect 373460 337588 373466 337652
rect 373993 337650 374059 337653
rect 374494 337650 374500 337652
rect 373993 337648 374500 337650
rect 373993 337592 373998 337648
rect 374054 337592 374500 337648
rect 373993 337590 374500 337592
rect 373993 337587 374059 337590
rect 374494 337588 374500 337590
rect 374564 337588 374570 337652
rect 376753 337650 376819 337653
rect 379513 337652 379579 337653
rect 376886 337650 376892 337652
rect 376753 337648 376892 337650
rect 376753 337592 376758 337648
rect 376814 337592 376892 337648
rect 376753 337590 376892 337592
rect 376753 337587 376819 337590
rect 376886 337588 376892 337590
rect 376956 337588 376962 337652
rect 379462 337588 379468 337652
rect 379532 337650 379579 337652
rect 380985 337650 381051 337653
rect 381118 337650 381124 337652
rect 379532 337648 379624 337650
rect 379574 337592 379624 337648
rect 379532 337590 379624 337592
rect 380985 337648 381124 337650
rect 380985 337592 380990 337648
rect 381046 337592 381124 337648
rect 380985 337590 381124 337592
rect 379532 337588 379579 337590
rect 379513 337587 379579 337588
rect 380985 337587 381051 337590
rect 381118 337588 381124 337590
rect 381188 337588 381194 337652
rect 383653 337650 383719 337653
rect 383878 337650 383884 337652
rect 383653 337648 383884 337650
rect 383653 337592 383658 337648
rect 383714 337592 383884 337648
rect 383653 337590 383884 337592
rect 383653 337587 383719 337590
rect 383878 337588 383884 337590
rect 383948 337588 383954 337652
rect 385033 337650 385099 337653
rect 385166 337650 385172 337652
rect 385033 337648 385172 337650
rect 385033 337592 385038 337648
rect 385094 337592 385172 337648
rect 385033 337590 385172 337592
rect 385033 337587 385099 337590
rect 385166 337588 385172 337590
rect 385236 337588 385242 337652
rect 386413 337650 386479 337653
rect 387558 337650 387564 337652
rect 386413 337648 387564 337650
rect 386413 337592 386418 337648
rect 386474 337592 387564 337648
rect 386413 337590 387564 337592
rect 386413 337587 386479 337590
rect 387558 337588 387564 337590
rect 387628 337588 387634 337652
rect 387885 337650 387951 337653
rect 388294 337650 388300 337652
rect 387885 337648 388300 337650
rect 387885 337592 387890 337648
rect 387946 337592 388300 337648
rect 387885 337590 388300 337592
rect 387885 337587 387951 337590
rect 388294 337588 388300 337590
rect 388364 337588 388370 337652
rect 389173 337650 389239 337653
rect 389766 337650 389772 337652
rect 389173 337648 389772 337650
rect 389173 337592 389178 337648
rect 389234 337592 389772 337648
rect 389173 337590 389772 337592
rect 389173 337587 389239 337590
rect 389766 337588 389772 337590
rect 389836 337588 389842 337652
rect 393405 337650 393471 337653
rect 393630 337650 393636 337652
rect 393405 337648 393636 337650
rect 393405 337592 393410 337648
rect 393466 337592 393636 337648
rect 393405 337590 393636 337592
rect 393405 337587 393471 337590
rect 393630 337588 393636 337590
rect 393700 337588 393706 337652
rect 396022 337588 396028 337652
rect 396092 337650 396098 337652
rect 396165 337650 396231 337653
rect 396092 337648 396231 337650
rect 396092 337592 396170 337648
rect 396226 337592 396231 337648
rect 396092 337590 396231 337592
rect 396092 337588 396098 337590
rect 396165 337587 396231 337590
rect 397545 337650 397611 337653
rect 398414 337650 398420 337652
rect 397545 337648 398420 337650
rect 397545 337592 397550 337648
rect 397606 337592 398420 337648
rect 397545 337590 398420 337592
rect 397545 337587 397611 337590
rect 398414 337588 398420 337590
rect 398484 337588 398490 337652
rect 402973 337650 403039 337653
rect 403566 337650 403572 337652
rect 402973 337648 403572 337650
rect 402973 337592 402978 337648
rect 403034 337592 403572 337648
rect 402973 337590 403572 337592
rect 402973 337587 403039 337590
rect 403566 337588 403572 337590
rect 403636 337588 403642 337652
rect 405733 337650 405799 337653
rect 405958 337650 405964 337652
rect 405733 337648 405964 337650
rect 405733 337592 405738 337648
rect 405794 337592 405964 337648
rect 405733 337590 405964 337592
rect 405733 337587 405799 337590
rect 405958 337588 405964 337590
rect 406028 337588 406034 337652
rect 409873 337650 409939 337653
rect 410926 337650 410932 337652
rect 409873 337648 410932 337650
rect 409873 337592 409878 337648
rect 409934 337592 410932 337648
rect 409873 337590 410932 337592
rect 409873 337587 409939 337590
rect 410926 337588 410932 337590
rect 410996 337588 411002 337652
rect 412633 337650 412699 337653
rect 413318 337650 413324 337652
rect 412633 337648 413324 337650
rect 412633 337592 412638 337648
rect 412694 337592 413324 337648
rect 412633 337590 413324 337592
rect 412633 337587 412699 337590
rect 413318 337588 413324 337590
rect 413388 337588 413394 337652
rect 415393 337650 415459 337653
rect 415894 337650 415900 337652
rect 415393 337648 415900 337650
rect 415393 337592 415398 337648
rect 415454 337592 415900 337648
rect 415393 337590 415900 337592
rect 415393 337587 415459 337590
rect 415894 337588 415900 337590
rect 415964 337588 415970 337652
rect 417417 337650 417483 337653
rect 420913 337652 420979 337653
rect 418286 337650 418292 337652
rect 417417 337648 418292 337650
rect 417417 337592 417422 337648
rect 417478 337592 418292 337648
rect 417417 337590 418292 337592
rect 417417 337587 417483 337590
rect 418286 337588 418292 337590
rect 418356 337588 418362 337652
rect 420862 337588 420868 337652
rect 420932 337650 420979 337652
rect 424317 337650 424383 337653
rect 425646 337650 425652 337652
rect 420932 337648 421024 337650
rect 420974 337592 421024 337648
rect 420932 337590 421024 337592
rect 424317 337648 425652 337650
rect 424317 337592 424322 337648
rect 424378 337592 425652 337648
rect 424317 337590 425652 337592
rect 420932 337588 420979 337590
rect 420913 337587 420979 337588
rect 424317 337587 424383 337590
rect 425646 337588 425652 337590
rect 425716 337588 425722 337652
rect 427813 337650 427879 337653
rect 428590 337650 428596 337652
rect 427813 337648 428596 337650
rect 427813 337592 427818 337648
rect 427874 337592 428596 337648
rect 427813 337590 428596 337592
rect 427813 337587 427879 337590
rect 428590 337588 428596 337590
rect 428660 337588 428666 337652
rect 430573 337650 430639 337653
rect 430982 337650 430988 337652
rect 430573 337648 430988 337650
rect 430573 337592 430578 337648
rect 430634 337592 430988 337648
rect 430573 337590 430988 337592
rect 430573 337587 430639 337590
rect 430982 337588 430988 337590
rect 431052 337588 431058 337652
rect 433333 337650 433399 337653
rect 433558 337650 433564 337652
rect 433333 337648 433564 337650
rect 433333 337592 433338 337648
rect 433394 337592 433564 337648
rect 433333 337590 433564 337592
rect 433333 337587 433399 337590
rect 433558 337588 433564 337590
rect 433628 337588 433634 337652
rect 440233 337650 440299 337653
rect 440918 337650 440924 337652
rect 440233 337648 440924 337650
rect 440233 337592 440238 337648
rect 440294 337592 440924 337648
rect 440233 337590 440924 337592
rect 440233 337587 440299 337590
rect 440918 337588 440924 337590
rect 440988 337588 440994 337652
rect 442993 337650 443059 337653
rect 443310 337650 443316 337652
rect 442993 337648 443316 337650
rect 442993 337592 442998 337648
rect 443054 337592 443316 337648
rect 442993 337590 443316 337592
rect 442993 337587 443059 337590
rect 443310 337588 443316 337590
rect 443380 337588 443386 337652
rect 57094 337452 57100 337516
rect 57164 337514 57170 337516
rect 57881 337514 57947 337517
rect 57164 337512 57947 337514
rect 57164 337456 57886 337512
rect 57942 337456 57947 337512
rect 57164 337454 57947 337456
rect 57164 337452 57170 337454
rect 57881 337451 57947 337454
rect 64270 337452 64276 337516
rect 64340 337514 64346 337516
rect 64781 337514 64847 337517
rect 64340 337512 64847 337514
rect 64340 337456 64786 337512
rect 64842 337456 64847 337512
rect 64340 337454 64847 337456
rect 64340 337452 64346 337454
rect 64781 337451 64847 337454
rect 72366 337452 72372 337516
rect 72436 337514 72442 337516
rect 72969 337514 73035 337517
rect 72436 337512 73035 337514
rect 72436 337456 72974 337512
rect 73030 337456 73035 337512
rect 72436 337454 73035 337456
rect 72436 337452 72442 337454
rect 72969 337451 73035 337454
rect 390553 337514 390619 337517
rect 390870 337514 390876 337516
rect 390553 337512 390876 337514
rect 390553 337456 390558 337512
rect 390614 337456 390876 337512
rect 390553 337454 390876 337456
rect 390553 337451 390619 337454
rect 390870 337452 390876 337454
rect 390940 337452 390946 337516
rect 393865 337514 393931 337517
rect 394366 337514 394372 337516
rect 393865 337512 394372 337514
rect 393865 337456 393870 337512
rect 393926 337456 394372 337512
rect 393865 337454 394372 337456
rect 393865 337451 393931 337454
rect 394366 337452 394372 337454
rect 394436 337452 394442 337516
rect 59445 337378 59511 337381
rect 60590 337378 60596 337380
rect 59445 337376 60596 337378
rect 59445 337320 59450 337376
rect 59506 337320 60596 337376
rect 59445 337318 60596 337320
rect 59445 337315 59511 337318
rect 60590 337316 60596 337318
rect 60660 337316 60666 337380
rect 69105 337378 69171 337381
rect 69974 337378 69980 337380
rect 69105 337376 69980 337378
rect 69105 337320 69110 337376
rect 69166 337320 69980 337376
rect 69105 337318 69980 337320
rect 69105 337315 69171 337318
rect 69974 337316 69980 337318
rect 70044 337316 70050 337380
rect 85982 337316 85988 337380
rect 86052 337378 86058 337380
rect 237414 337378 237420 337380
rect 86052 337318 237420 337378
rect 86052 337316 86058 337318
rect 237414 337316 237420 337318
rect 237484 337316 237490 337380
rect 380893 337378 380959 337381
rect 381670 337378 381676 337380
rect 380893 337376 381676 337378
rect 380893 337320 380898 337376
rect 380954 337320 381676 337376
rect 380893 337318 381676 337320
rect 380893 337315 380959 337318
rect 381670 337316 381676 337318
rect 381740 337316 381746 337380
rect 397453 337378 397519 337381
rect 398046 337378 398052 337380
rect 397453 337376 398052 337378
rect 397453 337320 397458 337376
rect 397514 337320 398052 337376
rect 397453 337318 398052 337320
rect 397453 337315 397519 337318
rect 398046 337316 398052 337318
rect 398116 337316 398122 337380
rect 59353 337242 59419 337245
rect 59486 337242 59492 337244
rect 59353 337240 59492 337242
rect 59353 337184 59358 337240
rect 59414 337184 59492 337240
rect 59353 337182 59492 337184
rect 59353 337179 59419 337182
rect 59486 337180 59492 337182
rect 59556 337180 59562 337244
rect 115974 337180 115980 337244
rect 116044 337242 116050 337244
rect 117221 337242 117287 337245
rect 116044 337240 117287 337242
rect 116044 337184 117226 337240
rect 117282 337184 117287 337240
rect 116044 337182 117287 337184
rect 116044 337180 116050 337182
rect 117221 337179 117287 337182
rect 375373 337242 375439 337245
rect 375782 337242 375788 337244
rect 375373 337240 375788 337242
rect 375373 337184 375378 337240
rect 375434 337184 375788 337240
rect 375373 337182 375788 337184
rect 375373 337179 375439 337182
rect 375782 337180 375788 337182
rect 375852 337180 375858 337244
rect 382273 337242 382339 337245
rect 383510 337242 383516 337244
rect 382273 337240 383516 337242
rect 382273 337184 382278 337240
rect 382334 337184 383516 337240
rect 382273 337182 383516 337184
rect 382273 337179 382339 337182
rect 383510 337180 383516 337182
rect 383580 337180 383586 337244
rect 445753 337242 445819 337245
rect 445886 337242 445892 337244
rect 445753 337240 445892 337242
rect 445753 337184 445758 337240
rect 445814 337184 445892 337240
rect 445753 337182 445892 337184
rect 445753 337179 445819 337182
rect 445886 337180 445892 337182
rect 445956 337180 445962 337244
rect 361573 337106 361639 337109
rect 361798 337106 361804 337108
rect 361573 337104 361804 337106
rect 361573 337048 361578 337104
rect 361634 337048 361804 337104
rect 361573 337046 361804 337048
rect 361573 337043 361639 337046
rect 361798 337044 361804 337046
rect 361868 337044 361874 337108
rect 375465 337106 375531 337109
rect 375966 337106 375972 337108
rect 375465 337104 375972 337106
rect 375465 337048 375470 337104
rect 375526 337048 375972 337104
rect 375465 337046 375972 337048
rect 375465 337043 375531 337046
rect 375966 337044 375972 337046
rect 376036 337044 376042 337108
rect 385125 337106 385191 337109
rect 385902 337106 385908 337108
rect 385125 337104 385908 337106
rect 385125 337048 385130 337104
rect 385186 337048 385908 337104
rect 385125 337046 385908 337048
rect 385125 337043 385191 337046
rect 385902 337044 385908 337046
rect 385972 337044 385978 337108
rect 434713 337106 434779 337109
rect 435766 337106 435772 337108
rect 434713 337104 435772 337106
rect 434713 337048 434718 337104
rect 434774 337048 435772 337104
rect 434713 337046 435772 337048
rect 434713 337043 434779 337046
rect 435766 337044 435772 337046
rect 435836 337044 435842 337108
rect 437473 337106 437539 337109
rect 438342 337106 438348 337108
rect 437473 337104 438348 337106
rect 437473 337048 437478 337104
rect 437534 337048 438348 337104
rect 437473 337046 438348 337048
rect 437473 337043 437539 337046
rect 438342 337044 438348 337046
rect 438412 337044 438418 337108
rect 82997 336970 83063 336973
rect 83590 336970 83596 336972
rect 82997 336968 83596 336970
rect 82997 336912 83002 336968
rect 83058 336912 83596 336968
rect 82997 336910 83596 336912
rect 82997 336907 83063 336910
rect 83590 336908 83596 336910
rect 83660 336908 83666 336972
rect 369853 336970 369919 336973
rect 370078 336970 370084 336972
rect 369853 336968 370084 336970
rect 369853 336912 369858 336968
rect 369914 336912 370084 336968
rect 369853 336910 370084 336912
rect 369853 336907 369919 336910
rect 370078 336908 370084 336910
rect 370148 336908 370154 336972
rect 392577 336970 392643 336973
rect 393446 336970 393452 336972
rect 392577 336968 393452 336970
rect 392577 336912 392582 336968
rect 392638 336912 393452 336968
rect 392577 336910 393452 336912
rect 392577 336907 392643 336910
rect 393446 336908 393452 336910
rect 393516 336908 393522 336972
rect 76046 336772 76052 336836
rect 76116 336834 76122 336836
rect 77201 336834 77267 336837
rect 81249 336836 81315 336837
rect 76116 336832 77267 336834
rect 76116 336776 77206 336832
rect 77262 336776 77267 336832
rect 76116 336774 77267 336776
rect 76116 336772 76122 336774
rect 77201 336771 77267 336774
rect 81198 336772 81204 336836
rect 81268 336834 81315 336836
rect 81268 336832 81360 336834
rect 81310 336776 81360 336832
rect 81268 336774 81360 336776
rect 81268 336772 81315 336774
rect 96102 336772 96108 336836
rect 96172 336834 96178 336836
rect 96521 336834 96587 336837
rect 96172 336832 96587 336834
rect 96172 336776 96526 336832
rect 96582 336776 96587 336832
rect 96172 336774 96587 336776
rect 96172 336772 96178 336774
rect 81249 336771 81315 336772
rect 96521 336771 96587 336774
rect 98862 336772 98868 336836
rect 98932 336834 98938 336836
rect 99281 336834 99347 336837
rect 98932 336832 99347 336834
rect 98932 336776 99286 336832
rect 99342 336776 99347 336832
rect 98932 336774 99347 336776
rect 98932 336772 98938 336774
rect 99281 336771 99347 336774
rect 103462 336772 103468 336836
rect 103532 336834 103538 336836
rect 104801 336834 104867 336837
rect 103532 336832 104867 336834
rect 103532 336776 104806 336832
rect 104862 336776 104867 336832
rect 103532 336774 104867 336776
rect 103532 336772 103538 336774
rect 104801 336771 104867 336774
rect 369945 336834 370011 336837
rect 370630 336834 370636 336836
rect 369945 336832 370636 336834
rect 369945 336776 369950 336832
rect 370006 336776 370636 336832
rect 369945 336774 370636 336776
rect 369945 336771 370011 336774
rect 370630 336772 370636 336774
rect 370700 336772 370706 336836
rect 400213 336834 400279 336837
rect 401174 336834 401180 336836
rect 400213 336832 401180 336834
rect 400213 336776 400218 336832
rect 400274 336776 401180 336832
rect 400213 336774 401180 336776
rect 400213 336771 400279 336774
rect 401174 336772 401180 336774
rect 401244 336772 401250 336836
rect 422661 336834 422727 336837
rect 423438 336834 423444 336836
rect 422661 336832 423444 336834
rect 422661 336776 422666 336832
rect 422722 336776 423444 336832
rect 422661 336774 423444 336776
rect 422661 336771 422727 336774
rect 423438 336772 423444 336774
rect 423508 336772 423514 336836
rect -960 332196 480 332436
rect 580165 325274 580231 325277
rect 583520 325274 584960 325364
rect 580165 325272 584960 325274
rect 580165 325216 580170 325272
rect 580226 325216 584960 325272
rect 580165 325214 584960 325216
rect 580165 325211 580231 325214
rect 583520 325124 584960 325214
rect -960 319290 480 319380
rect 3417 319290 3483 319293
rect -960 319288 3483 319290
rect -960 319232 3422 319288
rect 3478 319232 3483 319288
rect -960 319230 3483 319232
rect -960 319140 480 319230
rect 3417 319227 3483 319230
rect 580165 312082 580231 312085
rect 583520 312082 584960 312172
rect 580165 312080 584960 312082
rect 580165 312024 580170 312080
rect 580226 312024 584960 312080
rect 580165 312022 584960 312024
rect 580165 312019 580231 312022
rect 583520 311932 584960 312022
rect -960 306234 480 306324
rect 3417 306234 3483 306237
rect -960 306232 3483 306234
rect -960 306176 3422 306232
rect 3478 306176 3483 306232
rect -960 306174 3483 306176
rect -960 306084 480 306174
rect 3417 306171 3483 306174
rect 580165 298754 580231 298757
rect 583520 298754 584960 298844
rect 580165 298752 584960 298754
rect 580165 298696 580170 298752
rect 580226 298696 584960 298752
rect 580165 298694 584960 298696
rect 580165 298691 580231 298694
rect 583520 298604 584960 298694
rect -960 293178 480 293268
rect 3417 293178 3483 293181
rect -960 293176 3483 293178
rect -960 293120 3422 293176
rect 3478 293120 3483 293176
rect -960 293118 3483 293120
rect -960 293028 480 293118
rect 3417 293115 3483 293118
rect 583520 285276 584960 285516
rect -960 279972 480 280212
rect 579797 272234 579863 272237
rect 583520 272234 584960 272324
rect 579797 272232 584960 272234
rect 579797 272176 579802 272232
rect 579858 272176 584960 272232
rect 579797 272174 584960 272176
rect 579797 272171 579863 272174
rect 583520 272084 584960 272174
rect -960 267202 480 267292
rect 3049 267202 3115 267205
rect -960 267200 3115 267202
rect -960 267144 3054 267200
rect 3110 267144 3115 267200
rect -960 267142 3115 267144
rect -960 267052 480 267142
rect 3049 267139 3115 267142
rect 580165 258906 580231 258909
rect 583520 258906 584960 258996
rect 580165 258904 584960 258906
rect 580165 258848 580170 258904
rect 580226 258848 584960 258904
rect 580165 258846 584960 258848
rect 580165 258843 580231 258846
rect 583520 258756 584960 258846
rect -960 254146 480 254236
rect 3417 254146 3483 254149
rect -960 254144 3483 254146
rect -960 254088 3422 254144
rect 3478 254088 3483 254144
rect -960 254086 3483 254088
rect -960 253996 480 254086
rect 3417 254083 3483 254086
rect 579797 245578 579863 245581
rect 583520 245578 584960 245668
rect 579797 245576 584960 245578
rect 579797 245520 579802 245576
rect 579858 245520 584960 245576
rect 579797 245518 584960 245520
rect 579797 245515 579863 245518
rect 583520 245428 584960 245518
rect 41781 244354 41847 244357
rect 266997 244354 267063 244357
rect 41781 244352 267063 244354
rect 41781 244296 41786 244352
rect 41842 244296 267002 244352
rect 267058 244296 267063 244352
rect 41781 244294 267063 244296
rect 41781 244291 41847 244294
rect 266997 244291 267063 244294
rect 42558 242932 42564 242996
rect 42628 242994 42634 242996
rect 184841 242994 184907 242997
rect 42628 242992 184907 242994
rect 42628 242936 184846 242992
rect 184902 242936 184907 242992
rect 42628 242934 184907 242936
rect 42628 242932 42634 242934
rect 184841 242931 184907 242934
rect -960 241090 480 241180
rect 3417 241090 3483 241093
rect -960 241088 3483 241090
rect -960 241032 3422 241088
rect 3478 241032 3483 241088
rect -960 241030 3483 241032
rect -960 240940 480 241030
rect 3417 241027 3483 241030
rect 39941 239866 40007 239869
rect 39941 239864 40234 239866
rect 39941 239808 39946 239864
rect 40002 239808 40234 239864
rect 39941 239806 40234 239808
rect 39941 239803 40007 239806
rect 40174 239292 40234 239806
rect 239765 238914 239831 238917
rect 239292 238912 239831 238914
rect 239292 238856 239770 238912
rect 239826 238856 239831 238912
rect 239292 238854 239831 238856
rect 239765 238851 239831 238854
rect 37089 234970 37155 234973
rect 37089 234968 40204 234970
rect 37089 234912 37094 234968
rect 37150 234912 40204 234968
rect 37089 234910 40204 234912
rect 37089 234907 37155 234910
rect 242801 233610 242867 233613
rect 239292 233608 242867 233610
rect 239292 233552 242806 233608
rect 242862 233552 242867 233608
rect 239292 233550 242867 233552
rect 242801 233547 242867 233550
rect 579797 232386 579863 232389
rect 583520 232386 584960 232476
rect 579797 232384 584960 232386
rect 579797 232328 579802 232384
rect 579858 232328 584960 232384
rect 579797 232326 584960 232328
rect 579797 232323 579863 232326
rect 583520 232236 584960 232326
rect 39205 230618 39271 230621
rect 39205 230616 40204 230618
rect 39205 230560 39210 230616
rect 39266 230560 40204 230616
rect 39205 230558 40204 230560
rect 39205 230555 39271 230558
rect 240685 228306 240751 228309
rect 239292 228304 240751 228306
rect 239292 228248 240690 228304
rect 240746 228248 240751 228304
rect 239292 228246 240751 228248
rect 240685 228243 240751 228246
rect -960 227884 480 228124
rect 37181 226266 37247 226269
rect 37181 226264 40204 226266
rect 37181 226208 37186 226264
rect 37242 226208 40204 226264
rect 37181 226206 40204 226208
rect 37181 226203 37247 226206
rect 242801 223002 242867 223005
rect 239292 223000 242867 223002
rect 239292 222944 242806 223000
rect 242862 222944 242867 223000
rect 239292 222942 242867 222944
rect 242801 222939 242867 222942
rect 37825 221778 37891 221781
rect 37825 221776 40204 221778
rect 37825 221720 37830 221776
rect 37886 221720 40204 221776
rect 37825 221718 40204 221720
rect 37825 221715 37891 221718
rect 580441 219058 580507 219061
rect 583520 219058 584960 219148
rect 580441 219056 584960 219058
rect 580441 219000 580446 219056
rect 580502 219000 584960 219056
rect 580441 218998 584960 219000
rect 580441 218995 580507 218998
rect 583520 218908 584960 218998
rect 242801 217698 242867 217701
rect 239292 217696 242867 217698
rect 239292 217640 242806 217696
rect 242862 217640 242867 217696
rect 239292 217638 242867 217640
rect 242801 217635 242867 217638
rect 38009 217426 38075 217429
rect 38009 217424 40204 217426
rect 38009 217368 38014 217424
rect 38070 217368 40204 217424
rect 38009 217366 40204 217368
rect 38009 217363 38075 217366
rect -960 214978 480 215068
rect 3325 214978 3391 214981
rect -960 214976 3391 214978
rect -960 214920 3330 214976
rect 3386 214920 3391 214976
rect -960 214918 3391 214920
rect -960 214828 480 214918
rect 3325 214915 3391 214918
rect 36629 213074 36695 213077
rect 36629 213072 40204 213074
rect 36629 213016 36634 213072
rect 36690 213016 40204 213072
rect 36629 213014 40204 213016
rect 36629 213011 36695 213014
rect 241973 212394 242039 212397
rect 239292 212392 242039 212394
rect 239292 212336 241978 212392
rect 242034 212336 242039 212392
rect 239292 212334 242039 212336
rect 241973 212331 242039 212334
rect 39113 208722 39179 208725
rect 39113 208720 40204 208722
rect 39113 208664 39118 208720
rect 39174 208664 40204 208720
rect 39113 208662 40204 208664
rect 39113 208659 39179 208662
rect 242525 207090 242591 207093
rect 239292 207088 242591 207090
rect 239292 207032 242530 207088
rect 242586 207032 242591 207088
rect 239292 207030 242591 207032
rect 242525 207027 242591 207030
rect 579889 205730 579955 205733
rect 583520 205730 584960 205820
rect 579889 205728 584960 205730
rect 579889 205672 579894 205728
rect 579950 205672 584960 205728
rect 579889 205670 584960 205672
rect 579889 205667 579955 205670
rect 583520 205580 584960 205670
rect 39021 204370 39087 204373
rect 39021 204368 40204 204370
rect 39021 204312 39026 204368
rect 39082 204312 40204 204368
rect 39021 204310 40204 204312
rect 39021 204307 39087 204310
rect -960 201922 480 202012
rect 3417 201922 3483 201925
rect -960 201920 3483 201922
rect -960 201864 3422 201920
rect 3478 201864 3483 201920
rect -960 201862 3483 201864
rect -960 201772 480 201862
rect 3417 201859 3483 201862
rect 242433 201786 242499 201789
rect 239292 201784 242499 201786
rect 239292 201728 242438 201784
rect 242494 201728 242499 201784
rect 239292 201726 242499 201728
rect 242433 201723 242499 201726
rect 36721 199882 36787 199885
rect 36721 199880 40204 199882
rect 36721 199824 36726 199880
rect 36782 199824 40204 199880
rect 36721 199822 40204 199824
rect 36721 199819 36787 199822
rect 242341 196482 242407 196485
rect 239292 196480 242407 196482
rect 239292 196424 242346 196480
rect 242402 196424 242407 196480
rect 239292 196422 242407 196424
rect 242341 196419 242407 196422
rect 38009 195530 38075 195533
rect 38009 195528 40204 195530
rect 38009 195472 38014 195528
rect 38070 195472 40204 195528
rect 38009 195470 40204 195472
rect 38009 195467 38075 195470
rect 580165 192538 580231 192541
rect 583520 192538 584960 192628
rect 580165 192536 584960 192538
rect 580165 192480 580170 192536
rect 580226 192480 584960 192536
rect 580165 192478 584960 192480
rect 580165 192475 580231 192478
rect 583520 192388 584960 192478
rect 38009 191178 38075 191181
rect 241881 191178 241947 191181
rect 38009 191176 40204 191178
rect 38009 191120 38014 191176
rect 38070 191120 40204 191176
rect 38009 191118 40204 191120
rect 239292 191176 241947 191178
rect 239292 191120 241886 191176
rect 241942 191120 241947 191176
rect 239292 191118 241947 191120
rect 38009 191115 38075 191118
rect 241881 191115 241947 191118
rect -960 188866 480 188956
rect 3417 188866 3483 188869
rect -960 188864 3483 188866
rect -960 188808 3422 188864
rect 3478 188808 3483 188864
rect -960 188806 3483 188808
rect -960 188716 480 188806
rect 3417 188803 3483 188806
rect 37365 186826 37431 186829
rect 37365 186824 40204 186826
rect 37365 186768 37370 186824
rect 37426 186768 40204 186824
rect 37365 186766 40204 186768
rect 37365 186763 37431 186766
rect 242801 185874 242867 185877
rect 239292 185872 242867 185874
rect 239292 185816 242806 185872
rect 242862 185816 242867 185872
rect 239292 185814 242867 185816
rect 242801 185811 242867 185814
rect 38929 182338 38995 182341
rect 38929 182336 40204 182338
rect 38929 182280 38934 182336
rect 38990 182280 40204 182336
rect 38929 182278 40204 182280
rect 38929 182275 38995 182278
rect 242801 180570 242867 180573
rect 239292 180568 242867 180570
rect 239292 180512 242806 180568
rect 242862 180512 242867 180568
rect 239292 180510 242867 180512
rect 242801 180507 242867 180510
rect 580349 179210 580415 179213
rect 583520 179210 584960 179300
rect 580349 179208 584960 179210
rect 580349 179152 580354 179208
rect 580410 179152 584960 179208
rect 580349 179150 584960 179152
rect 580349 179147 580415 179150
rect 583520 179060 584960 179150
rect 38009 177986 38075 177989
rect 38009 177984 40204 177986
rect 38009 177928 38014 177984
rect 38070 177928 40204 177984
rect 38009 177926 40204 177928
rect 38009 177923 38075 177926
rect -960 175796 480 176036
rect 242801 175266 242867 175269
rect 239292 175264 242867 175266
rect 239292 175208 242806 175264
rect 242862 175208 242867 175264
rect 239292 175206 242867 175208
rect 242801 175203 242867 175206
rect 38009 173634 38075 173637
rect 38009 173632 40204 173634
rect 38009 173576 38014 173632
rect 38070 173576 40204 173632
rect 38009 173574 40204 173576
rect 38009 173571 38075 173574
rect 241881 169962 241947 169965
rect 239292 169960 241947 169962
rect 239292 169904 241886 169960
rect 241942 169904 241947 169960
rect 239292 169902 241947 169904
rect 241881 169899 241947 169902
rect 38009 169282 38075 169285
rect 38009 169280 40204 169282
rect 38009 169224 38014 169280
rect 38070 169224 40204 169280
rect 38009 169222 40204 169224
rect 38009 169219 38075 169222
rect 580165 165882 580231 165885
rect 583520 165882 584960 165972
rect 580165 165880 584960 165882
rect 580165 165824 580170 165880
rect 580226 165824 584960 165880
rect 580165 165822 584960 165824
rect 580165 165819 580231 165822
rect 583520 165732 584960 165822
rect 36813 164930 36879 164933
rect 36813 164928 40204 164930
rect 36813 164872 36818 164928
rect 36874 164872 40204 164928
rect 36813 164870 40204 164872
rect 36813 164867 36879 164870
rect 240593 164658 240659 164661
rect 239292 164656 240659 164658
rect 239292 164600 240598 164656
rect 240654 164600 240659 164656
rect 239292 164598 240659 164600
rect 240593 164595 240659 164598
rect -960 162890 480 162980
rect 3233 162890 3299 162893
rect -960 162888 3299 162890
rect -960 162832 3238 162888
rect 3294 162832 3299 162888
rect -960 162830 3299 162832
rect -960 162740 480 162830
rect 3233 162827 3299 162830
rect 38009 160442 38075 160445
rect 38009 160440 40204 160442
rect 38009 160384 38014 160440
rect 38070 160384 40204 160440
rect 38009 160382 40204 160384
rect 38009 160379 38075 160382
rect 241881 159354 241947 159357
rect 239292 159352 241947 159354
rect 239292 159296 241886 159352
rect 241942 159296 241947 159352
rect 239292 159294 241947 159296
rect 241881 159291 241947 159294
rect 36905 156090 36971 156093
rect 36905 156088 40204 156090
rect 36905 156032 36910 156088
rect 36966 156032 40204 156088
rect 36905 156030 40204 156032
rect 36905 156027 36971 156030
rect 240501 154050 240567 154053
rect 239292 154048 240567 154050
rect 239292 153992 240506 154048
rect 240562 153992 240567 154048
rect 239292 153990 240567 153992
rect 240501 153987 240567 153990
rect 579797 152690 579863 152693
rect 583520 152690 584960 152780
rect 579797 152688 584960 152690
rect 579797 152632 579802 152688
rect 579858 152632 584960 152688
rect 579797 152630 584960 152632
rect 579797 152627 579863 152630
rect 583520 152540 584960 152630
rect 38009 151738 38075 151741
rect 38009 151736 40204 151738
rect 38009 151680 38014 151736
rect 38070 151680 40204 151736
rect 38009 151678 40204 151680
rect 38009 151675 38075 151678
rect -960 149834 480 149924
rect 3417 149834 3483 149837
rect -960 149832 3483 149834
rect -960 149776 3422 149832
rect 3478 149776 3483 149832
rect -960 149774 3483 149776
rect -960 149684 480 149774
rect 3417 149771 3483 149774
rect 242801 148746 242867 148749
rect 239292 148744 242867 148746
rect 239292 148688 242806 148744
rect 242862 148688 242867 148744
rect 239292 148686 242867 148688
rect 242801 148683 242867 148686
rect 38009 147386 38075 147389
rect 38009 147384 40204 147386
rect 38009 147328 38014 147384
rect 38070 147328 40204 147384
rect 38009 147326 40204 147328
rect 38009 147323 38075 147326
rect 241881 143442 241947 143445
rect 239292 143440 241947 143442
rect 239292 143384 241886 143440
rect 241942 143384 241947 143440
rect 239292 143382 241947 143384
rect 241881 143379 241947 143382
rect 36997 143034 37063 143037
rect 36997 143032 40204 143034
rect 36997 142976 37002 143032
rect 37058 142976 40204 143032
rect 36997 142974 40204 142976
rect 36997 142971 37063 142974
rect 580165 139362 580231 139365
rect 583520 139362 584960 139452
rect 580165 139360 584960 139362
rect 580165 139304 580170 139360
rect 580226 139304 584960 139360
rect 580165 139302 584960 139304
rect 580165 139299 580231 139302
rect 583520 139212 584960 139302
rect 38009 138546 38075 138549
rect 38009 138544 40204 138546
rect 38009 138488 38014 138544
rect 38070 138488 40204 138544
rect 38009 138486 40204 138488
rect 38009 138483 38075 138486
rect 240409 138138 240475 138141
rect 239292 138136 240475 138138
rect 239292 138080 240414 138136
rect 240470 138080 240475 138136
rect 239292 138078 240475 138080
rect 240409 138075 240475 138078
rect -960 136778 480 136868
rect 3233 136778 3299 136781
rect -960 136776 3299 136778
rect -960 136720 3238 136776
rect 3294 136720 3299 136776
rect -960 136718 3299 136720
rect -960 136628 480 136718
rect 3233 136715 3299 136718
rect 38101 134194 38167 134197
rect 38101 134192 40204 134194
rect 38101 134136 38106 134192
rect 38162 134136 40204 134192
rect 38101 134134 40204 134136
rect 38101 134131 38167 134134
rect 243077 132834 243143 132837
rect 239292 132832 243143 132834
rect 239292 132776 243082 132832
rect 243138 132776 243143 132832
rect 239292 132774 243143 132776
rect 243077 132771 243143 132774
rect 38009 129842 38075 129845
rect 38009 129840 40204 129842
rect 38009 129784 38014 129840
rect 38070 129784 40204 129840
rect 38009 129782 40204 129784
rect 38009 129779 38075 129782
rect 242249 127530 242315 127533
rect 239292 127528 242315 127530
rect 239292 127472 242254 127528
rect 242310 127472 242315 127528
rect 239292 127470 242315 127472
rect 242249 127467 242315 127470
rect 580165 126034 580231 126037
rect 583520 126034 584960 126124
rect 580165 126032 584960 126034
rect 580165 125976 580170 126032
rect 580226 125976 584960 126032
rect 580165 125974 584960 125976
rect 580165 125971 580231 125974
rect 583520 125884 584960 125974
rect 38009 125490 38075 125493
rect 38009 125488 40204 125490
rect 38009 125432 38014 125488
rect 38070 125432 40204 125488
rect 38009 125430 40204 125432
rect 38009 125427 38075 125430
rect -960 123572 480 123812
rect 241973 122226 242039 122229
rect 239292 122224 242039 122226
rect 239292 122168 241978 122224
rect 242034 122168 242039 122224
rect 239292 122166 242039 122168
rect 241973 122163 242039 122166
rect 37917 121002 37983 121005
rect 37917 121000 40204 121002
rect 37917 120944 37922 121000
rect 37978 120944 40204 121000
rect 37917 120942 40204 120944
rect 37917 120939 37983 120942
rect 242801 116922 242867 116925
rect 239292 116920 242867 116922
rect 239292 116864 242806 116920
rect 242862 116864 242867 116920
rect 239292 116862 242867 116864
rect 242801 116859 242867 116862
rect 37733 116650 37799 116653
rect 37733 116648 40204 116650
rect 37733 116592 37738 116648
rect 37794 116592 40204 116648
rect 37733 116590 40204 116592
rect 37733 116587 37799 116590
rect 580165 112842 580231 112845
rect 583520 112842 584960 112932
rect 580165 112840 584960 112842
rect 580165 112784 580170 112840
rect 580226 112784 584960 112840
rect 580165 112782 584960 112784
rect 580165 112779 580231 112782
rect 583520 112692 584960 112782
rect 38009 112298 38075 112301
rect 38009 112296 40204 112298
rect 38009 112240 38014 112296
rect 38070 112240 40204 112296
rect 38009 112238 40204 112240
rect 38009 112235 38075 112238
rect 241881 111618 241947 111621
rect 239292 111616 241947 111618
rect 239292 111560 241886 111616
rect 241942 111560 241947 111616
rect 239292 111558 241947 111560
rect 241881 111555 241947 111558
rect -960 110666 480 110756
rect 3417 110666 3483 110669
rect -960 110664 3483 110666
rect -960 110608 3422 110664
rect 3478 110608 3483 110664
rect -960 110606 3483 110608
rect -960 110516 480 110606
rect 3417 110603 3483 110606
rect 37641 107946 37707 107949
rect 37641 107944 40204 107946
rect 37641 107888 37646 107944
rect 37702 107888 40204 107944
rect 37641 107886 40204 107888
rect 37641 107883 37707 107886
rect 241881 106314 241947 106317
rect 239292 106312 241947 106314
rect 239292 106256 241886 106312
rect 241942 106256 241947 106312
rect 239292 106254 241947 106256
rect 241881 106251 241947 106254
rect 38653 103594 38719 103597
rect 38653 103592 40204 103594
rect 38653 103536 38658 103592
rect 38714 103536 40204 103592
rect 38653 103534 40204 103536
rect 38653 103531 38719 103534
rect 241789 101010 241855 101013
rect 239292 101008 241855 101010
rect 239292 100952 241794 101008
rect 241850 100952 241855 101008
rect 239292 100950 241855 100952
rect 241789 100947 241855 100950
rect 580165 99514 580231 99517
rect 583520 99514 584960 99604
rect 580165 99512 584960 99514
rect 580165 99456 580170 99512
rect 580226 99456 584960 99512
rect 580165 99454 584960 99456
rect 580165 99451 580231 99454
rect 583520 99364 584960 99454
rect 38285 99106 38351 99109
rect 38285 99104 40204 99106
rect 38285 99048 38290 99104
rect 38346 99048 40204 99104
rect 38285 99046 40204 99048
rect 38285 99043 38351 99046
rect -960 97610 480 97700
rect 3417 97610 3483 97613
rect -960 97608 3483 97610
rect -960 97552 3422 97608
rect 3478 97552 3483 97608
rect -960 97550 3483 97552
rect -960 97460 480 97550
rect 3417 97547 3483 97550
rect 242801 95706 242867 95709
rect 239292 95704 242867 95706
rect 239292 95648 242806 95704
rect 242862 95648 242867 95704
rect 239292 95646 242867 95648
rect 242801 95643 242867 95646
rect 38009 94754 38075 94757
rect 38009 94752 40204 94754
rect 38009 94696 38014 94752
rect 38070 94696 40204 94752
rect 38009 94694 40204 94696
rect 38009 94691 38075 94694
rect 38009 90402 38075 90405
rect 242801 90402 242867 90405
rect 38009 90400 40204 90402
rect 38009 90344 38014 90400
rect 38070 90344 40204 90400
rect 38009 90342 40204 90344
rect 239292 90400 242867 90402
rect 239292 90344 242806 90400
rect 242862 90344 242867 90400
rect 239292 90342 242867 90344
rect 38009 90339 38075 90342
rect 242801 90339 242867 90342
rect 580165 86186 580231 86189
rect 583520 86186 584960 86276
rect 580165 86184 584960 86186
rect 580165 86128 580170 86184
rect 580226 86128 584960 86184
rect 580165 86126 584960 86128
rect 580165 86123 580231 86126
rect 38561 86050 38627 86053
rect 38561 86048 40204 86050
rect 38561 85992 38566 86048
rect 38622 85992 40204 86048
rect 583520 86036 584960 86126
rect 38561 85990 40204 85992
rect 38561 85987 38627 85990
rect 241513 85098 241579 85101
rect 239292 85096 241579 85098
rect 239292 85040 241518 85096
rect 241574 85040 241579 85096
rect 239292 85038 241579 85040
rect 241513 85035 241579 85038
rect -960 84690 480 84780
rect 3141 84690 3207 84693
rect -960 84688 3207 84690
rect -960 84632 3146 84688
rect 3202 84632 3207 84688
rect -960 84630 3207 84632
rect -960 84540 480 84630
rect 3141 84627 3207 84630
rect 38837 81562 38903 81565
rect 38837 81560 40204 81562
rect 38837 81504 38842 81560
rect 38898 81504 40204 81560
rect 38837 81502 40204 81504
rect 38837 81499 38903 81502
rect 242249 79794 242315 79797
rect 239292 79792 242315 79794
rect 239292 79736 242254 79792
rect 242310 79736 242315 79792
rect 239292 79734 242315 79736
rect 242249 79731 242315 79734
rect 38009 77210 38075 77213
rect 38009 77208 40204 77210
rect 38009 77152 38014 77208
rect 38070 77152 40204 77208
rect 38009 77150 40204 77152
rect 38009 77147 38075 77150
rect 241513 74490 241579 74493
rect 239292 74488 241579 74490
rect 239292 74432 241518 74488
rect 241574 74432 241579 74488
rect 239292 74430 241579 74432
rect 241513 74427 241579 74430
rect 579981 72994 580047 72997
rect 583520 72994 584960 73084
rect 579981 72992 584960 72994
rect 579981 72936 579986 72992
rect 580042 72936 584960 72992
rect 579981 72934 584960 72936
rect 579981 72931 580047 72934
rect 38745 72858 38811 72861
rect 38745 72856 40204 72858
rect 38745 72800 38750 72856
rect 38806 72800 40204 72856
rect 583520 72844 584960 72934
rect 38745 72798 40204 72800
rect 38745 72795 38811 72798
rect -960 71634 480 71724
rect 3417 71634 3483 71637
rect -960 71632 3483 71634
rect -960 71576 3422 71632
rect 3478 71576 3483 71632
rect -960 71574 3483 71576
rect -960 71484 480 71574
rect 3417 71571 3483 71574
rect 241697 69186 241763 69189
rect 239292 69184 241763 69186
rect 239292 69128 241702 69184
rect 241758 69128 241763 69184
rect 239292 69126 241763 69128
rect 241697 69123 241763 69126
rect 38009 68506 38075 68509
rect 38009 68504 40204 68506
rect 38009 68448 38014 68504
rect 38070 68448 40204 68504
rect 38009 68446 40204 68448
rect 38009 68443 38075 68446
rect 38193 64154 38259 64157
rect 38193 64152 40204 64154
rect 38193 64096 38198 64152
rect 38254 64096 40204 64152
rect 38193 64094 40204 64096
rect 38193 64091 38259 64094
rect 242801 63882 242867 63885
rect 239292 63880 242867 63882
rect 239292 63824 242806 63880
rect 242862 63824 242867 63880
rect 239292 63822 242867 63824
rect 242801 63819 242867 63822
rect 38009 59666 38075 59669
rect 580257 59666 580323 59669
rect 583520 59666 584960 59756
rect 38009 59664 40204 59666
rect 38009 59608 38014 59664
rect 38070 59608 40204 59664
rect 38009 59606 40204 59608
rect 580257 59664 584960 59666
rect 580257 59608 580262 59664
rect 580318 59608 584960 59664
rect 580257 59606 584960 59608
rect 38009 59603 38075 59606
rect 580257 59603 580323 59606
rect 583520 59516 584960 59606
rect -960 58578 480 58668
rect 3049 58578 3115 58581
rect 241513 58578 241579 58581
rect -960 58576 3115 58578
rect -960 58520 3054 58576
rect 3110 58520 3115 58576
rect -960 58518 3115 58520
rect 239292 58576 241579 58578
rect 239292 58520 241518 58576
rect 241574 58520 241579 58576
rect 239292 58518 241579 58520
rect -960 58428 480 58518
rect 3049 58515 3115 58518
rect 241513 58515 241579 58518
rect 38009 55314 38075 55317
rect 38009 55312 40204 55314
rect 38009 55256 38014 55312
rect 38070 55256 40204 55312
rect 38009 55254 40204 55256
rect 38009 55251 38075 55254
rect 241973 53274 242039 53277
rect 239292 53272 242039 53274
rect 239292 53216 241978 53272
rect 242034 53216 242039 53272
rect 239292 53214 242039 53216
rect 241973 53211 242039 53214
rect 37825 50962 37891 50965
rect 37825 50960 40204 50962
rect 37825 50904 37830 50960
rect 37886 50904 40204 50960
rect 37825 50902 40204 50904
rect 37825 50899 37891 50902
rect 241605 47970 241671 47973
rect 239292 47968 241671 47970
rect 239292 47912 241610 47968
rect 241666 47912 241671 47968
rect 239292 47910 241671 47912
rect 241605 47907 241671 47910
rect 38009 46610 38075 46613
rect 38009 46608 40204 46610
rect 38009 46552 38014 46608
rect 38070 46552 40204 46608
rect 38009 46550 40204 46552
rect 38009 46547 38075 46550
rect 580165 46338 580231 46341
rect 583520 46338 584960 46428
rect 580165 46336 584960 46338
rect 580165 46280 580170 46336
rect 580226 46280 584960 46336
rect 580165 46278 584960 46280
rect 580165 46275 580231 46278
rect 583520 46188 584960 46278
rect -960 45522 480 45612
rect 3417 45522 3483 45525
rect -960 45520 3483 45522
rect -960 45464 3422 45520
rect 3478 45464 3483 45520
rect -960 45462 3483 45464
rect -960 45372 480 45462
rect 3417 45459 3483 45462
rect 240317 42666 240383 42669
rect 239292 42664 240383 42666
rect 239292 42608 240322 42664
rect 240378 42608 240383 42664
rect 239292 42606 240383 42608
rect 240317 42603 240383 42606
rect 38009 42258 38075 42261
rect 38009 42256 40204 42258
rect 38009 42200 38014 42256
rect 38070 42200 40204 42256
rect 38009 42198 40204 42200
rect 38009 42195 38075 42198
rect 42057 39946 42123 39949
rect 42558 39946 42564 39948
rect 42057 39944 42564 39946
rect 42057 39888 42062 39944
rect 42118 39888 42564 39944
rect 42057 39886 42564 39888
rect 42057 39883 42123 39886
rect 42558 39884 42564 39886
rect 42628 39884 42634 39948
rect 41454 38524 41460 38588
rect 41524 38586 41530 38588
rect 42057 38586 42123 38589
rect 41524 38584 42123 38586
rect 41524 38528 42062 38584
rect 42118 38528 42123 38584
rect 41524 38526 42123 38528
rect 41524 38524 41530 38526
rect 42057 38523 42123 38526
rect 47710 38524 47716 38588
rect 47780 38586 47786 38588
rect 198733 38586 198799 38589
rect 47780 38584 198799 38586
rect 47780 38528 198738 38584
rect 198794 38528 198799 38584
rect 47780 38526 198799 38528
rect 47780 38524 47786 38526
rect 198733 38523 198799 38526
rect 235809 38586 235875 38589
rect 370497 38586 370563 38589
rect 235809 38584 370563 38586
rect 235809 38528 235814 38584
rect 235870 38528 370502 38584
rect 370558 38528 370563 38584
rect 235809 38526 370563 38528
rect 235809 38523 235875 38526
rect 370497 38523 370563 38526
rect 210141 38450 210207 38453
rect 237414 38450 237420 38452
rect 210141 38448 237420 38450
rect 210141 38392 210146 38448
rect 210202 38392 237420 38448
rect 210141 38390 237420 38392
rect 210141 38387 210207 38390
rect 237414 38388 237420 38390
rect 237484 38388 237490 38452
rect 580165 33146 580231 33149
rect 583520 33146 584960 33236
rect 580165 33144 584960 33146
rect 580165 33088 580170 33144
rect 580226 33088 584960 33144
rect 580165 33086 584960 33088
rect 580165 33083 580231 33086
rect 583520 32996 584960 33086
rect -960 32466 480 32556
rect 2773 32466 2839 32469
rect -960 32464 2839 32466
rect -960 32408 2778 32464
rect 2834 32408 2839 32464
rect -960 32406 2839 32408
rect -960 32316 480 32406
rect 2773 32403 2839 32406
rect 580165 19818 580231 19821
rect 583520 19818 584960 19908
rect 580165 19816 584960 19818
rect 580165 19760 580170 19816
rect 580226 19760 584960 19816
rect 580165 19758 584960 19760
rect 580165 19755 580231 19758
rect 583520 19668 584960 19758
rect -960 19410 480 19500
rect 3417 19410 3483 19413
rect -960 19408 3483 19410
rect -960 19352 3422 19408
rect 3478 19352 3483 19408
rect -960 19350 3483 19352
rect -960 19260 480 19350
rect 3417 19347 3483 19350
rect 580257 6626 580323 6629
rect 583520 6626 584960 6716
rect 580257 6624 584960 6626
rect -960 6490 480 6580
rect 580257 6568 580262 6624
rect 580318 6568 584960 6624
rect 580257 6566 584960 6568
rect 580257 6563 580323 6566
rect 3417 6490 3483 6493
rect -960 6488 3483 6490
rect -960 6432 3422 6488
rect 3478 6432 3483 6488
rect 583520 6476 584960 6566
rect -960 6430 3483 6432
rect -960 6340 480 6430
rect 3417 6427 3483 6430
rect 10317 6218 10383 6221
rect 41454 6218 41460 6220
rect 10317 6216 41460 6218
rect 10317 6160 10322 6216
rect 10378 6160 41460 6216
rect 10317 6158 41460 6160
rect 10317 6155 10383 6158
rect 41454 6156 41460 6158
rect 41524 6156 41530 6220
<< via3 >>
rect 76972 338132 77036 338196
rect 90956 338132 91020 338196
rect 131068 338132 131132 338196
rect 372292 338132 372356 338196
rect 382780 338132 382844 338196
rect 386460 338132 386524 338196
rect 408172 338132 408236 338196
rect 356100 338056 356164 338060
rect 356100 338000 356114 338056
rect 356114 338000 356164 338056
rect 356100 337996 356164 338000
rect 368980 337996 369044 338060
rect 55996 337860 56060 337924
rect 47716 337724 47780 337788
rect 68324 337860 68388 337924
rect 78076 337860 78140 337924
rect 97948 337860 98012 337924
rect 378548 337860 378612 337924
rect 392164 337860 392228 337924
rect 395660 337860 395724 337924
rect 396580 337860 396644 337924
rect 399156 337860 399220 337924
rect 67588 337724 67652 337788
rect 71268 337724 71332 337788
rect 73476 337724 73540 337788
rect 75868 337724 75932 337788
rect 82860 337724 82924 337788
rect 87644 337724 87708 337788
rect 91508 337724 91572 337788
rect 93348 337724 93412 337788
rect 94268 337724 94332 337788
rect 99052 337724 99116 337788
rect 143396 337724 143460 337788
rect 364196 337724 364260 337788
rect 368060 337724 368124 337788
rect 373580 337724 373644 337788
rect 377996 337724 378060 337788
rect 380572 337724 380636 337788
rect 388668 337724 388732 337788
rect 391060 337724 391124 337788
rect 58204 337588 58268 337652
rect 61884 337588 61948 337652
rect 63172 337588 63236 337652
rect 65380 337588 65444 337652
rect 66668 337588 66732 337652
rect 68692 337588 68756 337652
rect 70716 337588 70780 337652
rect 73660 337588 73724 337652
rect 74580 337588 74644 337652
rect 78444 337648 78508 337652
rect 78444 337592 78494 337648
rect 78494 337592 78508 337648
rect 78444 337588 78508 337592
rect 79548 337588 79612 337652
rect 81020 337648 81084 337652
rect 81020 337592 81070 337648
rect 81070 337592 81084 337648
rect 81020 337588 81084 337592
rect 81756 337588 81820 337652
rect 83412 337588 83476 337652
rect 85252 337648 85316 337652
rect 85252 337592 85302 337648
rect 85302 337592 85316 337648
rect 85252 337588 85316 337592
rect 86356 337648 86420 337652
rect 86356 337592 86406 337648
rect 86406 337592 86420 337648
rect 86356 337588 86420 337592
rect 88196 337648 88260 337652
rect 88196 337592 88210 337648
rect 88210 337592 88260 337648
rect 88196 337588 88260 337592
rect 88748 337588 88812 337652
rect 89852 337588 89916 337652
rect 92244 337588 92308 337652
rect 93532 337588 93596 337652
rect 95740 337588 95804 337652
rect 97028 337588 97092 337652
rect 100892 337588 100956 337652
rect 106044 337588 106108 337652
rect 108252 337588 108316 337652
rect 111012 337588 111076 337652
rect 113404 337588 113468 337652
rect 118556 337648 118620 337652
rect 118556 337592 118606 337648
rect 118606 337592 118620 337648
rect 118556 337588 118620 337592
rect 120948 337588 121012 337652
rect 123524 337588 123588 337652
rect 125916 337588 125980 337652
rect 128492 337588 128556 337652
rect 133460 337588 133524 337652
rect 135852 337588 135916 337652
rect 138612 337588 138676 337652
rect 141004 337588 141068 337652
rect 145972 337588 146036 337652
rect 357020 337588 357084 337652
rect 358124 337588 358188 337652
rect 359596 337588 359660 337652
rect 360516 337588 360580 337652
rect 363092 337588 363156 337652
rect 365484 337588 365548 337652
rect 366404 337588 366468 337652
rect 367508 337588 367572 337652
rect 371372 337648 371436 337652
rect 371372 337592 371386 337648
rect 371386 337592 371436 337648
rect 371372 337588 371436 337592
rect 373396 337588 373460 337652
rect 374500 337588 374564 337652
rect 376892 337588 376956 337652
rect 379468 337648 379532 337652
rect 379468 337592 379518 337648
rect 379518 337592 379532 337648
rect 379468 337588 379532 337592
rect 381124 337588 381188 337652
rect 383884 337588 383948 337652
rect 385172 337588 385236 337652
rect 387564 337588 387628 337652
rect 388300 337588 388364 337652
rect 389772 337588 389836 337652
rect 393636 337588 393700 337652
rect 396028 337588 396092 337652
rect 398420 337588 398484 337652
rect 403572 337588 403636 337652
rect 405964 337588 406028 337652
rect 410932 337588 410996 337652
rect 413324 337588 413388 337652
rect 415900 337588 415964 337652
rect 418292 337588 418356 337652
rect 420868 337648 420932 337652
rect 420868 337592 420918 337648
rect 420918 337592 420932 337648
rect 420868 337588 420932 337592
rect 425652 337588 425716 337652
rect 428596 337588 428660 337652
rect 430988 337588 431052 337652
rect 433564 337588 433628 337652
rect 440924 337588 440988 337652
rect 443316 337588 443380 337652
rect 57100 337452 57164 337516
rect 64276 337452 64340 337516
rect 72372 337452 72436 337516
rect 390876 337452 390940 337516
rect 394372 337452 394436 337516
rect 60596 337316 60660 337380
rect 69980 337316 70044 337380
rect 85988 337316 86052 337380
rect 237420 337316 237484 337380
rect 381676 337316 381740 337380
rect 398052 337316 398116 337380
rect 59492 337180 59556 337244
rect 115980 337180 116044 337244
rect 375788 337180 375852 337244
rect 383516 337180 383580 337244
rect 445892 337180 445956 337244
rect 361804 337044 361868 337108
rect 375972 337044 376036 337108
rect 385908 337044 385972 337108
rect 435772 337044 435836 337108
rect 438348 337044 438412 337108
rect 83596 336908 83660 336972
rect 370084 336908 370148 336972
rect 393452 336908 393516 336972
rect 76052 336772 76116 336836
rect 81204 336832 81268 336836
rect 81204 336776 81254 336832
rect 81254 336776 81268 336832
rect 81204 336772 81268 336776
rect 96108 336772 96172 336836
rect 98868 336772 98932 336836
rect 103468 336772 103532 336836
rect 370636 336772 370700 336836
rect 401180 336772 401244 336836
rect 423444 336772 423508 336836
rect 42564 242932 42628 242996
rect 42564 39884 42628 39948
rect 41460 38524 41524 38588
rect 47716 38524 47780 38588
rect 237420 38388 237484 38452
rect 41460 6156 41524 6220
<< metal4 >>
rect -8726 711558 -8106 711590
rect -8726 711322 -8694 711558
rect -8458 711322 -8374 711558
rect -8138 711322 -8106 711558
rect -8726 711238 -8106 711322
rect -8726 711002 -8694 711238
rect -8458 711002 -8374 711238
rect -8138 711002 -8106 711238
rect -8726 679394 -8106 711002
rect -8726 679158 -8694 679394
rect -8458 679158 -8374 679394
rect -8138 679158 -8106 679394
rect -8726 643394 -8106 679158
rect -8726 643158 -8694 643394
rect -8458 643158 -8374 643394
rect -8138 643158 -8106 643394
rect -8726 607394 -8106 643158
rect -8726 607158 -8694 607394
rect -8458 607158 -8374 607394
rect -8138 607158 -8106 607394
rect -8726 571394 -8106 607158
rect -8726 571158 -8694 571394
rect -8458 571158 -8374 571394
rect -8138 571158 -8106 571394
rect -8726 535394 -8106 571158
rect -8726 535158 -8694 535394
rect -8458 535158 -8374 535394
rect -8138 535158 -8106 535394
rect -8726 499394 -8106 535158
rect -8726 499158 -8694 499394
rect -8458 499158 -8374 499394
rect -8138 499158 -8106 499394
rect -8726 463394 -8106 499158
rect -8726 463158 -8694 463394
rect -8458 463158 -8374 463394
rect -8138 463158 -8106 463394
rect -8726 427394 -8106 463158
rect -8726 427158 -8694 427394
rect -8458 427158 -8374 427394
rect -8138 427158 -8106 427394
rect -8726 391394 -8106 427158
rect -8726 391158 -8694 391394
rect -8458 391158 -8374 391394
rect -8138 391158 -8106 391394
rect -8726 355394 -8106 391158
rect -8726 355158 -8694 355394
rect -8458 355158 -8374 355394
rect -8138 355158 -8106 355394
rect -8726 319394 -8106 355158
rect -8726 319158 -8694 319394
rect -8458 319158 -8374 319394
rect -8138 319158 -8106 319394
rect -8726 283394 -8106 319158
rect -8726 283158 -8694 283394
rect -8458 283158 -8374 283394
rect -8138 283158 -8106 283394
rect -8726 247394 -8106 283158
rect -8726 247158 -8694 247394
rect -8458 247158 -8374 247394
rect -8138 247158 -8106 247394
rect -8726 211394 -8106 247158
rect -8726 211158 -8694 211394
rect -8458 211158 -8374 211394
rect -8138 211158 -8106 211394
rect -8726 175394 -8106 211158
rect -8726 175158 -8694 175394
rect -8458 175158 -8374 175394
rect -8138 175158 -8106 175394
rect -8726 139394 -8106 175158
rect -8726 139158 -8694 139394
rect -8458 139158 -8374 139394
rect -8138 139158 -8106 139394
rect -8726 103394 -8106 139158
rect -8726 103158 -8694 103394
rect -8458 103158 -8374 103394
rect -8138 103158 -8106 103394
rect -8726 67394 -8106 103158
rect -8726 67158 -8694 67394
rect -8458 67158 -8374 67394
rect -8138 67158 -8106 67394
rect -8726 31394 -8106 67158
rect -8726 31158 -8694 31394
rect -8458 31158 -8374 31394
rect -8138 31158 -8106 31394
rect -8726 -7066 -8106 31158
rect -7766 710598 -7146 710630
rect -7766 710362 -7734 710598
rect -7498 710362 -7414 710598
rect -7178 710362 -7146 710598
rect -7766 710278 -7146 710362
rect -7766 710042 -7734 710278
rect -7498 710042 -7414 710278
rect -7178 710042 -7146 710278
rect -7766 697394 -7146 710042
rect 11904 710598 12504 711590
rect 11904 710362 12086 710598
rect 12322 710362 12504 710598
rect 11904 710278 12504 710362
rect 11904 710042 12086 710278
rect 12322 710042 12504 710278
rect -7766 697158 -7734 697394
rect -7498 697158 -7414 697394
rect -7178 697158 -7146 697394
rect -7766 661394 -7146 697158
rect -7766 661158 -7734 661394
rect -7498 661158 -7414 661394
rect -7178 661158 -7146 661394
rect -7766 625394 -7146 661158
rect -7766 625158 -7734 625394
rect -7498 625158 -7414 625394
rect -7178 625158 -7146 625394
rect -7766 589394 -7146 625158
rect -7766 589158 -7734 589394
rect -7498 589158 -7414 589394
rect -7178 589158 -7146 589394
rect -7766 553394 -7146 589158
rect -7766 553158 -7734 553394
rect -7498 553158 -7414 553394
rect -7178 553158 -7146 553394
rect -7766 517394 -7146 553158
rect -7766 517158 -7734 517394
rect -7498 517158 -7414 517394
rect -7178 517158 -7146 517394
rect -7766 481394 -7146 517158
rect -7766 481158 -7734 481394
rect -7498 481158 -7414 481394
rect -7178 481158 -7146 481394
rect -7766 445394 -7146 481158
rect -7766 445158 -7734 445394
rect -7498 445158 -7414 445394
rect -7178 445158 -7146 445394
rect -7766 409394 -7146 445158
rect -7766 409158 -7734 409394
rect -7498 409158 -7414 409394
rect -7178 409158 -7146 409394
rect -7766 373394 -7146 409158
rect -7766 373158 -7734 373394
rect -7498 373158 -7414 373394
rect -7178 373158 -7146 373394
rect -7766 337394 -7146 373158
rect -7766 337158 -7734 337394
rect -7498 337158 -7414 337394
rect -7178 337158 -7146 337394
rect -7766 301394 -7146 337158
rect -7766 301158 -7734 301394
rect -7498 301158 -7414 301394
rect -7178 301158 -7146 301394
rect -7766 265394 -7146 301158
rect -7766 265158 -7734 265394
rect -7498 265158 -7414 265394
rect -7178 265158 -7146 265394
rect -7766 229394 -7146 265158
rect -7766 229158 -7734 229394
rect -7498 229158 -7414 229394
rect -7178 229158 -7146 229394
rect -7766 193394 -7146 229158
rect -7766 193158 -7734 193394
rect -7498 193158 -7414 193394
rect -7178 193158 -7146 193394
rect -7766 157394 -7146 193158
rect -7766 157158 -7734 157394
rect -7498 157158 -7414 157394
rect -7178 157158 -7146 157394
rect -7766 121394 -7146 157158
rect -7766 121158 -7734 121394
rect -7498 121158 -7414 121394
rect -7178 121158 -7146 121394
rect -7766 85394 -7146 121158
rect -7766 85158 -7734 85394
rect -7498 85158 -7414 85394
rect -7178 85158 -7146 85394
rect -7766 49394 -7146 85158
rect -7766 49158 -7734 49394
rect -7498 49158 -7414 49394
rect -7178 49158 -7146 49394
rect -7766 13394 -7146 49158
rect -7766 13158 -7734 13394
rect -7498 13158 -7414 13394
rect -7178 13158 -7146 13394
rect -7766 -6106 -7146 13158
rect -6806 709638 -6186 709670
rect -6806 709402 -6774 709638
rect -6538 709402 -6454 709638
rect -6218 709402 -6186 709638
rect -6806 709318 -6186 709402
rect -6806 709082 -6774 709318
rect -6538 709082 -6454 709318
rect -6218 709082 -6186 709318
rect -6806 675694 -6186 709082
rect -6806 675458 -6774 675694
rect -6538 675458 -6454 675694
rect -6218 675458 -6186 675694
rect -6806 639694 -6186 675458
rect -6806 639458 -6774 639694
rect -6538 639458 -6454 639694
rect -6218 639458 -6186 639694
rect -6806 603694 -6186 639458
rect -6806 603458 -6774 603694
rect -6538 603458 -6454 603694
rect -6218 603458 -6186 603694
rect -6806 567694 -6186 603458
rect -6806 567458 -6774 567694
rect -6538 567458 -6454 567694
rect -6218 567458 -6186 567694
rect -6806 531694 -6186 567458
rect -6806 531458 -6774 531694
rect -6538 531458 -6454 531694
rect -6218 531458 -6186 531694
rect -6806 495694 -6186 531458
rect -6806 495458 -6774 495694
rect -6538 495458 -6454 495694
rect -6218 495458 -6186 495694
rect -6806 459694 -6186 495458
rect -6806 459458 -6774 459694
rect -6538 459458 -6454 459694
rect -6218 459458 -6186 459694
rect -6806 423694 -6186 459458
rect -6806 423458 -6774 423694
rect -6538 423458 -6454 423694
rect -6218 423458 -6186 423694
rect -6806 387694 -6186 423458
rect -6806 387458 -6774 387694
rect -6538 387458 -6454 387694
rect -6218 387458 -6186 387694
rect -6806 351694 -6186 387458
rect -6806 351458 -6774 351694
rect -6538 351458 -6454 351694
rect -6218 351458 -6186 351694
rect -6806 315694 -6186 351458
rect -6806 315458 -6774 315694
rect -6538 315458 -6454 315694
rect -6218 315458 -6186 315694
rect -6806 279694 -6186 315458
rect -6806 279458 -6774 279694
rect -6538 279458 -6454 279694
rect -6218 279458 -6186 279694
rect -6806 243694 -6186 279458
rect -6806 243458 -6774 243694
rect -6538 243458 -6454 243694
rect -6218 243458 -6186 243694
rect -6806 207694 -6186 243458
rect -6806 207458 -6774 207694
rect -6538 207458 -6454 207694
rect -6218 207458 -6186 207694
rect -6806 171694 -6186 207458
rect -6806 171458 -6774 171694
rect -6538 171458 -6454 171694
rect -6218 171458 -6186 171694
rect -6806 135694 -6186 171458
rect -6806 135458 -6774 135694
rect -6538 135458 -6454 135694
rect -6218 135458 -6186 135694
rect -6806 99694 -6186 135458
rect -6806 99458 -6774 99694
rect -6538 99458 -6454 99694
rect -6218 99458 -6186 99694
rect -6806 63694 -6186 99458
rect -6806 63458 -6774 63694
rect -6538 63458 -6454 63694
rect -6218 63458 -6186 63694
rect -6806 27694 -6186 63458
rect -6806 27458 -6774 27694
rect -6538 27458 -6454 27694
rect -6218 27458 -6186 27694
rect -6806 -5146 -6186 27458
rect -5846 708678 -5226 708710
rect -5846 708442 -5814 708678
rect -5578 708442 -5494 708678
rect -5258 708442 -5226 708678
rect -5846 708358 -5226 708442
rect -5846 708122 -5814 708358
rect -5578 708122 -5494 708358
rect -5258 708122 -5226 708358
rect -5846 693694 -5226 708122
rect 8204 708678 8804 709670
rect 8204 708442 8386 708678
rect 8622 708442 8804 708678
rect 8204 708358 8804 708442
rect 8204 708122 8386 708358
rect 8622 708122 8804 708358
rect -5846 693458 -5814 693694
rect -5578 693458 -5494 693694
rect -5258 693458 -5226 693694
rect -5846 657694 -5226 693458
rect -5846 657458 -5814 657694
rect -5578 657458 -5494 657694
rect -5258 657458 -5226 657694
rect -5846 621694 -5226 657458
rect -5846 621458 -5814 621694
rect -5578 621458 -5494 621694
rect -5258 621458 -5226 621694
rect -5846 585694 -5226 621458
rect -5846 585458 -5814 585694
rect -5578 585458 -5494 585694
rect -5258 585458 -5226 585694
rect -5846 549694 -5226 585458
rect -5846 549458 -5814 549694
rect -5578 549458 -5494 549694
rect -5258 549458 -5226 549694
rect -5846 513694 -5226 549458
rect -5846 513458 -5814 513694
rect -5578 513458 -5494 513694
rect -5258 513458 -5226 513694
rect -5846 477694 -5226 513458
rect -5846 477458 -5814 477694
rect -5578 477458 -5494 477694
rect -5258 477458 -5226 477694
rect -5846 441694 -5226 477458
rect -5846 441458 -5814 441694
rect -5578 441458 -5494 441694
rect -5258 441458 -5226 441694
rect -5846 405694 -5226 441458
rect -5846 405458 -5814 405694
rect -5578 405458 -5494 405694
rect -5258 405458 -5226 405694
rect -5846 369694 -5226 405458
rect -5846 369458 -5814 369694
rect -5578 369458 -5494 369694
rect -5258 369458 -5226 369694
rect -5846 333694 -5226 369458
rect -5846 333458 -5814 333694
rect -5578 333458 -5494 333694
rect -5258 333458 -5226 333694
rect -5846 297694 -5226 333458
rect -5846 297458 -5814 297694
rect -5578 297458 -5494 297694
rect -5258 297458 -5226 297694
rect -5846 261694 -5226 297458
rect -5846 261458 -5814 261694
rect -5578 261458 -5494 261694
rect -5258 261458 -5226 261694
rect -5846 225694 -5226 261458
rect -5846 225458 -5814 225694
rect -5578 225458 -5494 225694
rect -5258 225458 -5226 225694
rect -5846 189694 -5226 225458
rect -5846 189458 -5814 189694
rect -5578 189458 -5494 189694
rect -5258 189458 -5226 189694
rect -5846 153694 -5226 189458
rect -5846 153458 -5814 153694
rect -5578 153458 -5494 153694
rect -5258 153458 -5226 153694
rect -5846 117694 -5226 153458
rect -5846 117458 -5814 117694
rect -5578 117458 -5494 117694
rect -5258 117458 -5226 117694
rect -5846 81694 -5226 117458
rect -5846 81458 -5814 81694
rect -5578 81458 -5494 81694
rect -5258 81458 -5226 81694
rect -5846 45694 -5226 81458
rect -5846 45458 -5814 45694
rect -5578 45458 -5494 45694
rect -5258 45458 -5226 45694
rect -5846 9694 -5226 45458
rect -5846 9458 -5814 9694
rect -5578 9458 -5494 9694
rect -5258 9458 -5226 9694
rect -5846 -4186 -5226 9458
rect -4886 707718 -4266 707750
rect -4886 707482 -4854 707718
rect -4618 707482 -4534 707718
rect -4298 707482 -4266 707718
rect -4886 707398 -4266 707482
rect -4886 707162 -4854 707398
rect -4618 707162 -4534 707398
rect -4298 707162 -4266 707398
rect -4886 671994 -4266 707162
rect -4886 671758 -4854 671994
rect -4618 671758 -4534 671994
rect -4298 671758 -4266 671994
rect -4886 635994 -4266 671758
rect -4886 635758 -4854 635994
rect -4618 635758 -4534 635994
rect -4298 635758 -4266 635994
rect -4886 599994 -4266 635758
rect -4886 599758 -4854 599994
rect -4618 599758 -4534 599994
rect -4298 599758 -4266 599994
rect -4886 563994 -4266 599758
rect -4886 563758 -4854 563994
rect -4618 563758 -4534 563994
rect -4298 563758 -4266 563994
rect -4886 527994 -4266 563758
rect -4886 527758 -4854 527994
rect -4618 527758 -4534 527994
rect -4298 527758 -4266 527994
rect -4886 491994 -4266 527758
rect -4886 491758 -4854 491994
rect -4618 491758 -4534 491994
rect -4298 491758 -4266 491994
rect -4886 455994 -4266 491758
rect -4886 455758 -4854 455994
rect -4618 455758 -4534 455994
rect -4298 455758 -4266 455994
rect -4886 419994 -4266 455758
rect -4886 419758 -4854 419994
rect -4618 419758 -4534 419994
rect -4298 419758 -4266 419994
rect -4886 383994 -4266 419758
rect -4886 383758 -4854 383994
rect -4618 383758 -4534 383994
rect -4298 383758 -4266 383994
rect -4886 347994 -4266 383758
rect -4886 347758 -4854 347994
rect -4618 347758 -4534 347994
rect -4298 347758 -4266 347994
rect -4886 311994 -4266 347758
rect -4886 311758 -4854 311994
rect -4618 311758 -4534 311994
rect -4298 311758 -4266 311994
rect -4886 275994 -4266 311758
rect -4886 275758 -4854 275994
rect -4618 275758 -4534 275994
rect -4298 275758 -4266 275994
rect -4886 239994 -4266 275758
rect -4886 239758 -4854 239994
rect -4618 239758 -4534 239994
rect -4298 239758 -4266 239994
rect -4886 203994 -4266 239758
rect -4886 203758 -4854 203994
rect -4618 203758 -4534 203994
rect -4298 203758 -4266 203994
rect -4886 167994 -4266 203758
rect -4886 167758 -4854 167994
rect -4618 167758 -4534 167994
rect -4298 167758 -4266 167994
rect -4886 131994 -4266 167758
rect -4886 131758 -4854 131994
rect -4618 131758 -4534 131994
rect -4298 131758 -4266 131994
rect -4886 95994 -4266 131758
rect -4886 95758 -4854 95994
rect -4618 95758 -4534 95994
rect -4298 95758 -4266 95994
rect -4886 59994 -4266 95758
rect -4886 59758 -4854 59994
rect -4618 59758 -4534 59994
rect -4298 59758 -4266 59994
rect -4886 23994 -4266 59758
rect -4886 23758 -4854 23994
rect -4618 23758 -4534 23994
rect -4298 23758 -4266 23994
rect -4886 -3226 -4266 23758
rect -3926 706758 -3306 706790
rect -3926 706522 -3894 706758
rect -3658 706522 -3574 706758
rect -3338 706522 -3306 706758
rect -3926 706438 -3306 706522
rect -3926 706202 -3894 706438
rect -3658 706202 -3574 706438
rect -3338 706202 -3306 706438
rect -3926 689994 -3306 706202
rect 4504 706758 5104 707750
rect 4504 706522 4686 706758
rect 4922 706522 5104 706758
rect 4504 706438 5104 706522
rect 4504 706202 4686 706438
rect 4922 706202 5104 706438
rect -3926 689758 -3894 689994
rect -3658 689758 -3574 689994
rect -3338 689758 -3306 689994
rect -3926 653994 -3306 689758
rect -3926 653758 -3894 653994
rect -3658 653758 -3574 653994
rect -3338 653758 -3306 653994
rect -3926 617994 -3306 653758
rect -3926 617758 -3894 617994
rect -3658 617758 -3574 617994
rect -3338 617758 -3306 617994
rect -3926 581994 -3306 617758
rect -3926 581758 -3894 581994
rect -3658 581758 -3574 581994
rect -3338 581758 -3306 581994
rect -3926 545994 -3306 581758
rect -3926 545758 -3894 545994
rect -3658 545758 -3574 545994
rect -3338 545758 -3306 545994
rect -3926 509994 -3306 545758
rect -3926 509758 -3894 509994
rect -3658 509758 -3574 509994
rect -3338 509758 -3306 509994
rect -3926 473994 -3306 509758
rect -3926 473758 -3894 473994
rect -3658 473758 -3574 473994
rect -3338 473758 -3306 473994
rect -3926 437994 -3306 473758
rect -3926 437758 -3894 437994
rect -3658 437758 -3574 437994
rect -3338 437758 -3306 437994
rect -3926 401994 -3306 437758
rect -3926 401758 -3894 401994
rect -3658 401758 -3574 401994
rect -3338 401758 -3306 401994
rect -3926 365994 -3306 401758
rect -3926 365758 -3894 365994
rect -3658 365758 -3574 365994
rect -3338 365758 -3306 365994
rect -3926 329994 -3306 365758
rect -3926 329758 -3894 329994
rect -3658 329758 -3574 329994
rect -3338 329758 -3306 329994
rect -3926 293994 -3306 329758
rect -3926 293758 -3894 293994
rect -3658 293758 -3574 293994
rect -3338 293758 -3306 293994
rect -3926 257994 -3306 293758
rect -3926 257758 -3894 257994
rect -3658 257758 -3574 257994
rect -3338 257758 -3306 257994
rect -3926 221994 -3306 257758
rect -3926 221758 -3894 221994
rect -3658 221758 -3574 221994
rect -3338 221758 -3306 221994
rect -3926 185994 -3306 221758
rect -3926 185758 -3894 185994
rect -3658 185758 -3574 185994
rect -3338 185758 -3306 185994
rect -3926 149994 -3306 185758
rect -3926 149758 -3894 149994
rect -3658 149758 -3574 149994
rect -3338 149758 -3306 149994
rect -3926 113994 -3306 149758
rect -3926 113758 -3894 113994
rect -3658 113758 -3574 113994
rect -3338 113758 -3306 113994
rect -3926 77994 -3306 113758
rect -3926 77758 -3894 77994
rect -3658 77758 -3574 77994
rect -3338 77758 -3306 77994
rect -3926 41994 -3306 77758
rect -3926 41758 -3894 41994
rect -3658 41758 -3574 41994
rect -3338 41758 -3306 41994
rect -3926 5994 -3306 41758
rect -3926 5758 -3894 5994
rect -3658 5758 -3574 5994
rect -3338 5758 -3306 5994
rect -3926 -2266 -3306 5758
rect -2966 705798 -2346 705830
rect -2966 705562 -2934 705798
rect -2698 705562 -2614 705798
rect -2378 705562 -2346 705798
rect -2966 705478 -2346 705562
rect -2966 705242 -2934 705478
rect -2698 705242 -2614 705478
rect -2378 705242 -2346 705478
rect -2966 668294 -2346 705242
rect -2966 668058 -2934 668294
rect -2698 668058 -2614 668294
rect -2378 668058 -2346 668294
rect -2966 632294 -2346 668058
rect -2966 632058 -2934 632294
rect -2698 632058 -2614 632294
rect -2378 632058 -2346 632294
rect -2966 596294 -2346 632058
rect -2966 596058 -2934 596294
rect -2698 596058 -2614 596294
rect -2378 596058 -2346 596294
rect -2966 560294 -2346 596058
rect -2966 560058 -2934 560294
rect -2698 560058 -2614 560294
rect -2378 560058 -2346 560294
rect -2966 524294 -2346 560058
rect -2966 524058 -2934 524294
rect -2698 524058 -2614 524294
rect -2378 524058 -2346 524294
rect -2966 488294 -2346 524058
rect -2966 488058 -2934 488294
rect -2698 488058 -2614 488294
rect -2378 488058 -2346 488294
rect -2966 452294 -2346 488058
rect -2966 452058 -2934 452294
rect -2698 452058 -2614 452294
rect -2378 452058 -2346 452294
rect -2966 416294 -2346 452058
rect -2966 416058 -2934 416294
rect -2698 416058 -2614 416294
rect -2378 416058 -2346 416294
rect -2966 380294 -2346 416058
rect -2966 380058 -2934 380294
rect -2698 380058 -2614 380294
rect -2378 380058 -2346 380294
rect -2966 344294 -2346 380058
rect -2966 344058 -2934 344294
rect -2698 344058 -2614 344294
rect -2378 344058 -2346 344294
rect -2966 308294 -2346 344058
rect -2966 308058 -2934 308294
rect -2698 308058 -2614 308294
rect -2378 308058 -2346 308294
rect -2966 272294 -2346 308058
rect -2966 272058 -2934 272294
rect -2698 272058 -2614 272294
rect -2378 272058 -2346 272294
rect -2966 236294 -2346 272058
rect -2966 236058 -2934 236294
rect -2698 236058 -2614 236294
rect -2378 236058 -2346 236294
rect -2966 200294 -2346 236058
rect -2966 200058 -2934 200294
rect -2698 200058 -2614 200294
rect -2378 200058 -2346 200294
rect -2966 164294 -2346 200058
rect -2966 164058 -2934 164294
rect -2698 164058 -2614 164294
rect -2378 164058 -2346 164294
rect -2966 128294 -2346 164058
rect -2966 128058 -2934 128294
rect -2698 128058 -2614 128294
rect -2378 128058 -2346 128294
rect -2966 92294 -2346 128058
rect -2966 92058 -2934 92294
rect -2698 92058 -2614 92294
rect -2378 92058 -2346 92294
rect -2966 56294 -2346 92058
rect -2966 56058 -2934 56294
rect -2698 56058 -2614 56294
rect -2378 56058 -2346 56294
rect -2966 20294 -2346 56058
rect -2966 20058 -2934 20294
rect -2698 20058 -2614 20294
rect -2378 20058 -2346 20294
rect -2966 -1306 -2346 20058
rect -2006 704838 -1386 704870
rect -2006 704602 -1974 704838
rect -1738 704602 -1654 704838
rect -1418 704602 -1386 704838
rect -2006 704518 -1386 704602
rect -2006 704282 -1974 704518
rect -1738 704282 -1654 704518
rect -1418 704282 -1386 704518
rect -2006 686294 -1386 704282
rect -2006 686058 -1974 686294
rect -1738 686058 -1654 686294
rect -1418 686058 -1386 686294
rect -2006 650294 -1386 686058
rect -2006 650058 -1974 650294
rect -1738 650058 -1654 650294
rect -1418 650058 -1386 650294
rect -2006 614294 -1386 650058
rect -2006 614058 -1974 614294
rect -1738 614058 -1654 614294
rect -1418 614058 -1386 614294
rect -2006 578294 -1386 614058
rect -2006 578058 -1974 578294
rect -1738 578058 -1654 578294
rect -1418 578058 -1386 578294
rect -2006 542294 -1386 578058
rect -2006 542058 -1974 542294
rect -1738 542058 -1654 542294
rect -1418 542058 -1386 542294
rect -2006 506294 -1386 542058
rect -2006 506058 -1974 506294
rect -1738 506058 -1654 506294
rect -1418 506058 -1386 506294
rect -2006 470294 -1386 506058
rect -2006 470058 -1974 470294
rect -1738 470058 -1654 470294
rect -1418 470058 -1386 470294
rect -2006 434294 -1386 470058
rect -2006 434058 -1974 434294
rect -1738 434058 -1654 434294
rect -1418 434058 -1386 434294
rect -2006 398294 -1386 434058
rect -2006 398058 -1974 398294
rect -1738 398058 -1654 398294
rect -1418 398058 -1386 398294
rect -2006 362294 -1386 398058
rect -2006 362058 -1974 362294
rect -1738 362058 -1654 362294
rect -1418 362058 -1386 362294
rect -2006 326294 -1386 362058
rect -2006 326058 -1974 326294
rect -1738 326058 -1654 326294
rect -1418 326058 -1386 326294
rect -2006 290294 -1386 326058
rect -2006 290058 -1974 290294
rect -1738 290058 -1654 290294
rect -1418 290058 -1386 290294
rect -2006 254294 -1386 290058
rect -2006 254058 -1974 254294
rect -1738 254058 -1654 254294
rect -1418 254058 -1386 254294
rect -2006 218294 -1386 254058
rect -2006 218058 -1974 218294
rect -1738 218058 -1654 218294
rect -1418 218058 -1386 218294
rect -2006 182294 -1386 218058
rect -2006 182058 -1974 182294
rect -1738 182058 -1654 182294
rect -1418 182058 -1386 182294
rect -2006 146294 -1386 182058
rect -2006 146058 -1974 146294
rect -1738 146058 -1654 146294
rect -1418 146058 -1386 146294
rect -2006 110294 -1386 146058
rect -2006 110058 -1974 110294
rect -1738 110058 -1654 110294
rect -1418 110058 -1386 110294
rect -2006 74294 -1386 110058
rect -2006 74058 -1974 74294
rect -1738 74058 -1654 74294
rect -1418 74058 -1386 74294
rect -2006 38294 -1386 74058
rect -2006 38058 -1974 38294
rect -1738 38058 -1654 38294
rect -1418 38058 -1386 38294
rect -2006 2294 -1386 38058
rect -2006 2058 -1974 2294
rect -1738 2058 -1654 2294
rect -1418 2058 -1386 2294
rect -2006 -346 -1386 2058
rect -2006 -582 -1974 -346
rect -1738 -582 -1654 -346
rect -1418 -582 -1386 -346
rect -2006 -666 -1386 -582
rect -2006 -902 -1974 -666
rect -1738 -902 -1654 -666
rect -1418 -902 -1386 -666
rect -2006 -934 -1386 -902
rect 804 704838 1404 705830
rect 804 704602 986 704838
rect 1222 704602 1404 704838
rect 804 704518 1404 704602
rect 804 704282 986 704518
rect 1222 704282 1404 704518
rect 804 686294 1404 704282
rect 804 686058 986 686294
rect 1222 686058 1404 686294
rect 804 650294 1404 686058
rect 804 650058 986 650294
rect 1222 650058 1404 650294
rect 804 614294 1404 650058
rect 804 614058 986 614294
rect 1222 614058 1404 614294
rect 804 578294 1404 614058
rect 804 578058 986 578294
rect 1222 578058 1404 578294
rect 804 542294 1404 578058
rect 804 542058 986 542294
rect 1222 542058 1404 542294
rect 804 506294 1404 542058
rect 804 506058 986 506294
rect 1222 506058 1404 506294
rect 804 470294 1404 506058
rect 804 470058 986 470294
rect 1222 470058 1404 470294
rect 804 434294 1404 470058
rect 804 434058 986 434294
rect 1222 434058 1404 434294
rect 804 398294 1404 434058
rect 804 398058 986 398294
rect 1222 398058 1404 398294
rect 804 362294 1404 398058
rect 804 362058 986 362294
rect 1222 362058 1404 362294
rect 804 326294 1404 362058
rect 804 326058 986 326294
rect 1222 326058 1404 326294
rect 804 290294 1404 326058
rect 804 290058 986 290294
rect 1222 290058 1404 290294
rect 804 254294 1404 290058
rect 804 254058 986 254294
rect 1222 254058 1404 254294
rect 804 218294 1404 254058
rect 804 218058 986 218294
rect 1222 218058 1404 218294
rect 804 182294 1404 218058
rect 804 182058 986 182294
rect 1222 182058 1404 182294
rect 804 146294 1404 182058
rect 804 146058 986 146294
rect 1222 146058 1404 146294
rect 804 110294 1404 146058
rect 804 110058 986 110294
rect 1222 110058 1404 110294
rect 804 74294 1404 110058
rect 804 74058 986 74294
rect 1222 74058 1404 74294
rect 804 38294 1404 74058
rect 804 38058 986 38294
rect 1222 38058 1404 38294
rect 804 2294 1404 38058
rect 804 2058 986 2294
rect 1222 2058 1404 2294
rect 804 -346 1404 2058
rect 804 -582 986 -346
rect 1222 -582 1404 -346
rect 804 -666 1404 -582
rect 804 -902 986 -666
rect 1222 -902 1404 -666
rect -2966 -1542 -2934 -1306
rect -2698 -1542 -2614 -1306
rect -2378 -1542 -2346 -1306
rect -2966 -1626 -2346 -1542
rect -2966 -1862 -2934 -1626
rect -2698 -1862 -2614 -1626
rect -2378 -1862 -2346 -1626
rect -2966 -1894 -2346 -1862
rect 804 -1894 1404 -902
rect 4504 689994 5104 706202
rect 4504 689758 4686 689994
rect 4922 689758 5104 689994
rect 4504 653994 5104 689758
rect 4504 653758 4686 653994
rect 4922 653758 5104 653994
rect 4504 617994 5104 653758
rect 4504 617758 4686 617994
rect 4922 617758 5104 617994
rect 4504 581994 5104 617758
rect 4504 581758 4686 581994
rect 4922 581758 5104 581994
rect 4504 545994 5104 581758
rect 4504 545758 4686 545994
rect 4922 545758 5104 545994
rect 4504 509994 5104 545758
rect 4504 509758 4686 509994
rect 4922 509758 5104 509994
rect 4504 473994 5104 509758
rect 4504 473758 4686 473994
rect 4922 473758 5104 473994
rect 4504 437994 5104 473758
rect 4504 437758 4686 437994
rect 4922 437758 5104 437994
rect 4504 401994 5104 437758
rect 4504 401758 4686 401994
rect 4922 401758 5104 401994
rect 4504 365994 5104 401758
rect 4504 365758 4686 365994
rect 4922 365758 5104 365994
rect 4504 329994 5104 365758
rect 4504 329758 4686 329994
rect 4922 329758 5104 329994
rect 4504 293994 5104 329758
rect 4504 293758 4686 293994
rect 4922 293758 5104 293994
rect 4504 257994 5104 293758
rect 4504 257758 4686 257994
rect 4922 257758 5104 257994
rect 4504 221994 5104 257758
rect 4504 221758 4686 221994
rect 4922 221758 5104 221994
rect 4504 185994 5104 221758
rect 4504 185758 4686 185994
rect 4922 185758 5104 185994
rect 4504 149994 5104 185758
rect 4504 149758 4686 149994
rect 4922 149758 5104 149994
rect 4504 113994 5104 149758
rect 4504 113758 4686 113994
rect 4922 113758 5104 113994
rect 4504 77994 5104 113758
rect 4504 77758 4686 77994
rect 4922 77758 5104 77994
rect 4504 41994 5104 77758
rect 4504 41758 4686 41994
rect 4922 41758 5104 41994
rect 4504 5994 5104 41758
rect 4504 5758 4686 5994
rect 4922 5758 5104 5994
rect -3926 -2502 -3894 -2266
rect -3658 -2502 -3574 -2266
rect -3338 -2502 -3306 -2266
rect -3926 -2586 -3306 -2502
rect -3926 -2822 -3894 -2586
rect -3658 -2822 -3574 -2586
rect -3338 -2822 -3306 -2586
rect -3926 -2854 -3306 -2822
rect 4504 -2266 5104 5758
rect 4504 -2502 4686 -2266
rect 4922 -2502 5104 -2266
rect 4504 -2586 5104 -2502
rect 4504 -2822 4686 -2586
rect 4922 -2822 5104 -2586
rect -4886 -3462 -4854 -3226
rect -4618 -3462 -4534 -3226
rect -4298 -3462 -4266 -3226
rect -4886 -3546 -4266 -3462
rect -4886 -3782 -4854 -3546
rect -4618 -3782 -4534 -3546
rect -4298 -3782 -4266 -3546
rect -4886 -3814 -4266 -3782
rect 4504 -3814 5104 -2822
rect 8204 693694 8804 708122
rect 8204 693458 8386 693694
rect 8622 693458 8804 693694
rect 8204 657694 8804 693458
rect 8204 657458 8386 657694
rect 8622 657458 8804 657694
rect 8204 621694 8804 657458
rect 8204 621458 8386 621694
rect 8622 621458 8804 621694
rect 8204 585694 8804 621458
rect 8204 585458 8386 585694
rect 8622 585458 8804 585694
rect 8204 549694 8804 585458
rect 8204 549458 8386 549694
rect 8622 549458 8804 549694
rect 8204 513694 8804 549458
rect 8204 513458 8386 513694
rect 8622 513458 8804 513694
rect 8204 477694 8804 513458
rect 8204 477458 8386 477694
rect 8622 477458 8804 477694
rect 8204 441694 8804 477458
rect 8204 441458 8386 441694
rect 8622 441458 8804 441694
rect 8204 405694 8804 441458
rect 8204 405458 8386 405694
rect 8622 405458 8804 405694
rect 8204 369694 8804 405458
rect 8204 369458 8386 369694
rect 8622 369458 8804 369694
rect 8204 333694 8804 369458
rect 8204 333458 8386 333694
rect 8622 333458 8804 333694
rect 8204 297694 8804 333458
rect 8204 297458 8386 297694
rect 8622 297458 8804 297694
rect 8204 261694 8804 297458
rect 8204 261458 8386 261694
rect 8622 261458 8804 261694
rect 8204 225694 8804 261458
rect 8204 225458 8386 225694
rect 8622 225458 8804 225694
rect 8204 189694 8804 225458
rect 8204 189458 8386 189694
rect 8622 189458 8804 189694
rect 8204 153694 8804 189458
rect 8204 153458 8386 153694
rect 8622 153458 8804 153694
rect 8204 117694 8804 153458
rect 8204 117458 8386 117694
rect 8622 117458 8804 117694
rect 8204 81694 8804 117458
rect 8204 81458 8386 81694
rect 8622 81458 8804 81694
rect 8204 45694 8804 81458
rect 8204 45458 8386 45694
rect 8622 45458 8804 45694
rect 8204 9694 8804 45458
rect 8204 9458 8386 9694
rect 8622 9458 8804 9694
rect -5846 -4422 -5814 -4186
rect -5578 -4422 -5494 -4186
rect -5258 -4422 -5226 -4186
rect -5846 -4506 -5226 -4422
rect -5846 -4742 -5814 -4506
rect -5578 -4742 -5494 -4506
rect -5258 -4742 -5226 -4506
rect -5846 -4774 -5226 -4742
rect 8204 -4186 8804 9458
rect 8204 -4422 8386 -4186
rect 8622 -4422 8804 -4186
rect 8204 -4506 8804 -4422
rect 8204 -4742 8386 -4506
rect 8622 -4742 8804 -4506
rect -6806 -5382 -6774 -5146
rect -6538 -5382 -6454 -5146
rect -6218 -5382 -6186 -5146
rect -6806 -5466 -6186 -5382
rect -6806 -5702 -6774 -5466
rect -6538 -5702 -6454 -5466
rect -6218 -5702 -6186 -5466
rect -6806 -5734 -6186 -5702
rect 8204 -5734 8804 -4742
rect 11904 697394 12504 710042
rect 29904 711558 30504 711590
rect 29904 711322 30086 711558
rect 30322 711322 30504 711558
rect 29904 711238 30504 711322
rect 29904 711002 30086 711238
rect 30322 711002 30504 711238
rect 26204 709638 26804 709670
rect 26204 709402 26386 709638
rect 26622 709402 26804 709638
rect 26204 709318 26804 709402
rect 26204 709082 26386 709318
rect 26622 709082 26804 709318
rect 22504 707718 23104 707750
rect 22504 707482 22686 707718
rect 22922 707482 23104 707718
rect 22504 707398 23104 707482
rect 22504 707162 22686 707398
rect 22922 707162 23104 707398
rect 11904 697158 12086 697394
rect 12322 697158 12504 697394
rect 11904 661394 12504 697158
rect 11904 661158 12086 661394
rect 12322 661158 12504 661394
rect 11904 625394 12504 661158
rect 11904 625158 12086 625394
rect 12322 625158 12504 625394
rect 11904 589394 12504 625158
rect 11904 589158 12086 589394
rect 12322 589158 12504 589394
rect 11904 553394 12504 589158
rect 11904 553158 12086 553394
rect 12322 553158 12504 553394
rect 11904 517394 12504 553158
rect 11904 517158 12086 517394
rect 12322 517158 12504 517394
rect 11904 481394 12504 517158
rect 11904 481158 12086 481394
rect 12322 481158 12504 481394
rect 11904 445394 12504 481158
rect 11904 445158 12086 445394
rect 12322 445158 12504 445394
rect 11904 409394 12504 445158
rect 11904 409158 12086 409394
rect 12322 409158 12504 409394
rect 11904 373394 12504 409158
rect 11904 373158 12086 373394
rect 12322 373158 12504 373394
rect 11904 337394 12504 373158
rect 11904 337158 12086 337394
rect 12322 337158 12504 337394
rect 11904 301394 12504 337158
rect 11904 301158 12086 301394
rect 12322 301158 12504 301394
rect 11904 265394 12504 301158
rect 11904 265158 12086 265394
rect 12322 265158 12504 265394
rect 11904 229394 12504 265158
rect 11904 229158 12086 229394
rect 12322 229158 12504 229394
rect 11904 193394 12504 229158
rect 11904 193158 12086 193394
rect 12322 193158 12504 193394
rect 11904 157394 12504 193158
rect 11904 157158 12086 157394
rect 12322 157158 12504 157394
rect 11904 121394 12504 157158
rect 11904 121158 12086 121394
rect 12322 121158 12504 121394
rect 11904 85394 12504 121158
rect 11904 85158 12086 85394
rect 12322 85158 12504 85394
rect 11904 49394 12504 85158
rect 11904 49158 12086 49394
rect 12322 49158 12504 49394
rect 11904 13394 12504 49158
rect 11904 13158 12086 13394
rect 12322 13158 12504 13394
rect -7766 -6342 -7734 -6106
rect -7498 -6342 -7414 -6106
rect -7178 -6342 -7146 -6106
rect -7766 -6426 -7146 -6342
rect -7766 -6662 -7734 -6426
rect -7498 -6662 -7414 -6426
rect -7178 -6662 -7146 -6426
rect -7766 -6694 -7146 -6662
rect 11904 -6106 12504 13158
rect 18804 705798 19404 705830
rect 18804 705562 18986 705798
rect 19222 705562 19404 705798
rect 18804 705478 19404 705562
rect 18804 705242 18986 705478
rect 19222 705242 19404 705478
rect 18804 668294 19404 705242
rect 18804 668058 18986 668294
rect 19222 668058 19404 668294
rect 18804 632294 19404 668058
rect 18804 632058 18986 632294
rect 19222 632058 19404 632294
rect 18804 596294 19404 632058
rect 18804 596058 18986 596294
rect 19222 596058 19404 596294
rect 18804 560294 19404 596058
rect 18804 560058 18986 560294
rect 19222 560058 19404 560294
rect 18804 524294 19404 560058
rect 18804 524058 18986 524294
rect 19222 524058 19404 524294
rect 18804 488294 19404 524058
rect 18804 488058 18986 488294
rect 19222 488058 19404 488294
rect 18804 452294 19404 488058
rect 18804 452058 18986 452294
rect 19222 452058 19404 452294
rect 18804 416294 19404 452058
rect 18804 416058 18986 416294
rect 19222 416058 19404 416294
rect 18804 380294 19404 416058
rect 18804 380058 18986 380294
rect 19222 380058 19404 380294
rect 18804 344294 19404 380058
rect 18804 344058 18986 344294
rect 19222 344058 19404 344294
rect 18804 308294 19404 344058
rect 18804 308058 18986 308294
rect 19222 308058 19404 308294
rect 18804 272294 19404 308058
rect 18804 272058 18986 272294
rect 19222 272058 19404 272294
rect 18804 236294 19404 272058
rect 18804 236058 18986 236294
rect 19222 236058 19404 236294
rect 18804 200294 19404 236058
rect 18804 200058 18986 200294
rect 19222 200058 19404 200294
rect 18804 164294 19404 200058
rect 18804 164058 18986 164294
rect 19222 164058 19404 164294
rect 18804 128294 19404 164058
rect 18804 128058 18986 128294
rect 19222 128058 19404 128294
rect 18804 92294 19404 128058
rect 18804 92058 18986 92294
rect 19222 92058 19404 92294
rect 18804 56294 19404 92058
rect 18804 56058 18986 56294
rect 19222 56058 19404 56294
rect 18804 20294 19404 56058
rect 18804 20058 18986 20294
rect 19222 20058 19404 20294
rect 18804 -1306 19404 20058
rect 18804 -1542 18986 -1306
rect 19222 -1542 19404 -1306
rect 18804 -1626 19404 -1542
rect 18804 -1862 18986 -1626
rect 19222 -1862 19404 -1626
rect 18804 -1894 19404 -1862
rect 22504 671994 23104 707162
rect 22504 671758 22686 671994
rect 22922 671758 23104 671994
rect 22504 635994 23104 671758
rect 22504 635758 22686 635994
rect 22922 635758 23104 635994
rect 22504 599994 23104 635758
rect 22504 599758 22686 599994
rect 22922 599758 23104 599994
rect 22504 563994 23104 599758
rect 22504 563758 22686 563994
rect 22922 563758 23104 563994
rect 22504 527994 23104 563758
rect 22504 527758 22686 527994
rect 22922 527758 23104 527994
rect 22504 491994 23104 527758
rect 22504 491758 22686 491994
rect 22922 491758 23104 491994
rect 22504 455994 23104 491758
rect 22504 455758 22686 455994
rect 22922 455758 23104 455994
rect 22504 419994 23104 455758
rect 22504 419758 22686 419994
rect 22922 419758 23104 419994
rect 22504 383994 23104 419758
rect 22504 383758 22686 383994
rect 22922 383758 23104 383994
rect 22504 347994 23104 383758
rect 22504 347758 22686 347994
rect 22922 347758 23104 347994
rect 22504 311994 23104 347758
rect 22504 311758 22686 311994
rect 22922 311758 23104 311994
rect 22504 275994 23104 311758
rect 22504 275758 22686 275994
rect 22922 275758 23104 275994
rect 22504 239994 23104 275758
rect 22504 239758 22686 239994
rect 22922 239758 23104 239994
rect 22504 203994 23104 239758
rect 22504 203758 22686 203994
rect 22922 203758 23104 203994
rect 22504 167994 23104 203758
rect 22504 167758 22686 167994
rect 22922 167758 23104 167994
rect 22504 131994 23104 167758
rect 22504 131758 22686 131994
rect 22922 131758 23104 131994
rect 22504 95994 23104 131758
rect 22504 95758 22686 95994
rect 22922 95758 23104 95994
rect 22504 59994 23104 95758
rect 22504 59758 22686 59994
rect 22922 59758 23104 59994
rect 22504 23994 23104 59758
rect 22504 23758 22686 23994
rect 22922 23758 23104 23994
rect 22504 -3226 23104 23758
rect 22504 -3462 22686 -3226
rect 22922 -3462 23104 -3226
rect 22504 -3546 23104 -3462
rect 22504 -3782 22686 -3546
rect 22922 -3782 23104 -3546
rect 22504 -3814 23104 -3782
rect 26204 675694 26804 709082
rect 26204 675458 26386 675694
rect 26622 675458 26804 675694
rect 26204 639694 26804 675458
rect 26204 639458 26386 639694
rect 26622 639458 26804 639694
rect 26204 603694 26804 639458
rect 26204 603458 26386 603694
rect 26622 603458 26804 603694
rect 26204 567694 26804 603458
rect 26204 567458 26386 567694
rect 26622 567458 26804 567694
rect 26204 531694 26804 567458
rect 26204 531458 26386 531694
rect 26622 531458 26804 531694
rect 26204 495694 26804 531458
rect 26204 495458 26386 495694
rect 26622 495458 26804 495694
rect 26204 459694 26804 495458
rect 26204 459458 26386 459694
rect 26622 459458 26804 459694
rect 26204 423694 26804 459458
rect 26204 423458 26386 423694
rect 26622 423458 26804 423694
rect 26204 387694 26804 423458
rect 26204 387458 26386 387694
rect 26622 387458 26804 387694
rect 26204 351694 26804 387458
rect 26204 351458 26386 351694
rect 26622 351458 26804 351694
rect 26204 315694 26804 351458
rect 26204 315458 26386 315694
rect 26622 315458 26804 315694
rect 26204 279694 26804 315458
rect 26204 279458 26386 279694
rect 26622 279458 26804 279694
rect 26204 243694 26804 279458
rect 26204 243458 26386 243694
rect 26622 243458 26804 243694
rect 26204 207694 26804 243458
rect 26204 207458 26386 207694
rect 26622 207458 26804 207694
rect 26204 171694 26804 207458
rect 26204 171458 26386 171694
rect 26622 171458 26804 171694
rect 26204 135694 26804 171458
rect 26204 135458 26386 135694
rect 26622 135458 26804 135694
rect 26204 99694 26804 135458
rect 26204 99458 26386 99694
rect 26622 99458 26804 99694
rect 26204 63694 26804 99458
rect 26204 63458 26386 63694
rect 26622 63458 26804 63694
rect 26204 27694 26804 63458
rect 26204 27458 26386 27694
rect 26622 27458 26804 27694
rect 26204 -5146 26804 27458
rect 26204 -5382 26386 -5146
rect 26622 -5382 26804 -5146
rect 26204 -5466 26804 -5382
rect 26204 -5702 26386 -5466
rect 26622 -5702 26804 -5466
rect 26204 -5734 26804 -5702
rect 29904 679394 30504 711002
rect 47904 710598 48504 711590
rect 47904 710362 48086 710598
rect 48322 710362 48504 710598
rect 47904 710278 48504 710362
rect 47904 710042 48086 710278
rect 48322 710042 48504 710278
rect 44204 708678 44804 709670
rect 44204 708442 44386 708678
rect 44622 708442 44804 708678
rect 44204 708358 44804 708442
rect 44204 708122 44386 708358
rect 44622 708122 44804 708358
rect 40504 706758 41104 707750
rect 40504 706522 40686 706758
rect 40922 706522 41104 706758
rect 40504 706438 41104 706522
rect 40504 706202 40686 706438
rect 40922 706202 41104 706438
rect 29904 679158 30086 679394
rect 30322 679158 30504 679394
rect 29904 643394 30504 679158
rect 29904 643158 30086 643394
rect 30322 643158 30504 643394
rect 29904 607394 30504 643158
rect 29904 607158 30086 607394
rect 30322 607158 30504 607394
rect 29904 571394 30504 607158
rect 29904 571158 30086 571394
rect 30322 571158 30504 571394
rect 29904 535394 30504 571158
rect 29904 535158 30086 535394
rect 30322 535158 30504 535394
rect 29904 499394 30504 535158
rect 29904 499158 30086 499394
rect 30322 499158 30504 499394
rect 29904 463394 30504 499158
rect 29904 463158 30086 463394
rect 30322 463158 30504 463394
rect 29904 427394 30504 463158
rect 29904 427158 30086 427394
rect 30322 427158 30504 427394
rect 29904 391394 30504 427158
rect 29904 391158 30086 391394
rect 30322 391158 30504 391394
rect 29904 355394 30504 391158
rect 29904 355158 30086 355394
rect 30322 355158 30504 355394
rect 29904 319394 30504 355158
rect 29904 319158 30086 319394
rect 30322 319158 30504 319394
rect 29904 283394 30504 319158
rect 29904 283158 30086 283394
rect 30322 283158 30504 283394
rect 29904 247394 30504 283158
rect 29904 247158 30086 247394
rect 30322 247158 30504 247394
rect 29904 211394 30504 247158
rect 29904 211158 30086 211394
rect 30322 211158 30504 211394
rect 29904 175394 30504 211158
rect 29904 175158 30086 175394
rect 30322 175158 30504 175394
rect 29904 139394 30504 175158
rect 29904 139158 30086 139394
rect 30322 139158 30504 139394
rect 29904 103394 30504 139158
rect 29904 103158 30086 103394
rect 30322 103158 30504 103394
rect 29904 67394 30504 103158
rect 29904 67158 30086 67394
rect 30322 67158 30504 67394
rect 29904 31394 30504 67158
rect 29904 31158 30086 31394
rect 30322 31158 30504 31394
rect 11904 -6342 12086 -6106
rect 12322 -6342 12504 -6106
rect 11904 -6426 12504 -6342
rect 11904 -6662 12086 -6426
rect 12322 -6662 12504 -6426
rect -8726 -7302 -8694 -7066
rect -8458 -7302 -8374 -7066
rect -8138 -7302 -8106 -7066
rect -8726 -7386 -8106 -7302
rect -8726 -7622 -8694 -7386
rect -8458 -7622 -8374 -7386
rect -8138 -7622 -8106 -7386
rect -8726 -7654 -8106 -7622
rect 11904 -7654 12504 -6662
rect 29904 -7066 30504 31158
rect 36804 704838 37404 705830
rect 36804 704602 36986 704838
rect 37222 704602 37404 704838
rect 36804 704518 37404 704602
rect 36804 704282 36986 704518
rect 37222 704282 37404 704518
rect 36804 686294 37404 704282
rect 36804 686058 36986 686294
rect 37222 686058 37404 686294
rect 36804 650294 37404 686058
rect 36804 650058 36986 650294
rect 37222 650058 37404 650294
rect 36804 614294 37404 650058
rect 36804 614058 36986 614294
rect 37222 614058 37404 614294
rect 36804 578294 37404 614058
rect 36804 578058 36986 578294
rect 37222 578058 37404 578294
rect 36804 542294 37404 578058
rect 36804 542058 36986 542294
rect 37222 542058 37404 542294
rect 36804 506294 37404 542058
rect 36804 506058 36986 506294
rect 37222 506058 37404 506294
rect 36804 470294 37404 506058
rect 36804 470058 36986 470294
rect 37222 470058 37404 470294
rect 36804 434294 37404 470058
rect 36804 434058 36986 434294
rect 37222 434058 37404 434294
rect 36804 398294 37404 434058
rect 40504 689994 41104 706202
rect 40504 689758 40686 689994
rect 40922 689758 41104 689994
rect 40504 653994 41104 689758
rect 40504 653758 40686 653994
rect 40922 653758 41104 653994
rect 40504 617994 41104 653758
rect 40504 617758 40686 617994
rect 40922 617758 41104 617994
rect 40504 581994 41104 617758
rect 40504 581758 40686 581994
rect 40922 581758 41104 581994
rect 40504 545994 41104 581758
rect 40504 545758 40686 545994
rect 40922 545758 41104 545994
rect 40504 509994 41104 545758
rect 40504 509758 40686 509994
rect 40922 509758 41104 509994
rect 40504 473994 41104 509758
rect 40504 473758 40686 473994
rect 40922 473758 41104 473994
rect 40504 437994 41104 473758
rect 40504 437758 40686 437994
rect 40922 437758 41104 437994
rect 40504 425308 41104 437758
rect 44204 693694 44804 708122
rect 44204 693458 44386 693694
rect 44622 693458 44804 693694
rect 44204 657694 44804 693458
rect 44204 657458 44386 657694
rect 44622 657458 44804 657694
rect 44204 621694 44804 657458
rect 44204 621458 44386 621694
rect 44622 621458 44804 621694
rect 44204 585694 44804 621458
rect 44204 585458 44386 585694
rect 44622 585458 44804 585694
rect 44204 549694 44804 585458
rect 44204 549458 44386 549694
rect 44622 549458 44804 549694
rect 44204 513694 44804 549458
rect 44204 513458 44386 513694
rect 44622 513458 44804 513694
rect 44204 477694 44804 513458
rect 44204 477458 44386 477694
rect 44622 477458 44804 477694
rect 44204 441694 44804 477458
rect 44204 441458 44386 441694
rect 44622 441458 44804 441694
rect 44204 425308 44804 441458
rect 47904 697394 48504 710042
rect 65904 711558 66504 711590
rect 65904 711322 66086 711558
rect 66322 711322 66504 711558
rect 65904 711238 66504 711322
rect 65904 711002 66086 711238
rect 66322 711002 66504 711238
rect 62204 709638 62804 709670
rect 62204 709402 62386 709638
rect 62622 709402 62804 709638
rect 62204 709318 62804 709402
rect 62204 709082 62386 709318
rect 62622 709082 62804 709318
rect 58504 707718 59104 707750
rect 58504 707482 58686 707718
rect 58922 707482 59104 707718
rect 58504 707398 59104 707482
rect 58504 707162 58686 707398
rect 58922 707162 59104 707398
rect 47904 697158 48086 697394
rect 48322 697158 48504 697394
rect 47904 661394 48504 697158
rect 47904 661158 48086 661394
rect 48322 661158 48504 661394
rect 47904 625394 48504 661158
rect 47904 625158 48086 625394
rect 48322 625158 48504 625394
rect 47904 589394 48504 625158
rect 47904 589158 48086 589394
rect 48322 589158 48504 589394
rect 47904 553394 48504 589158
rect 47904 553158 48086 553394
rect 48322 553158 48504 553394
rect 47904 517394 48504 553158
rect 47904 517158 48086 517394
rect 48322 517158 48504 517394
rect 47904 481394 48504 517158
rect 47904 481158 48086 481394
rect 48322 481158 48504 481394
rect 47904 445394 48504 481158
rect 47904 445158 48086 445394
rect 48322 445158 48504 445394
rect 47904 425308 48504 445158
rect 54804 705798 55404 705830
rect 54804 705562 54986 705798
rect 55222 705562 55404 705798
rect 54804 705478 55404 705562
rect 54804 705242 54986 705478
rect 55222 705242 55404 705478
rect 54804 668294 55404 705242
rect 54804 668058 54986 668294
rect 55222 668058 55404 668294
rect 54804 632294 55404 668058
rect 54804 632058 54986 632294
rect 55222 632058 55404 632294
rect 54804 596294 55404 632058
rect 54804 596058 54986 596294
rect 55222 596058 55404 596294
rect 54804 560294 55404 596058
rect 54804 560058 54986 560294
rect 55222 560058 55404 560294
rect 54804 524294 55404 560058
rect 54804 524058 54986 524294
rect 55222 524058 55404 524294
rect 54804 488294 55404 524058
rect 54804 488058 54986 488294
rect 55222 488058 55404 488294
rect 54804 452294 55404 488058
rect 54804 452058 54986 452294
rect 55222 452058 55404 452294
rect 54804 425308 55404 452058
rect 58504 671994 59104 707162
rect 58504 671758 58686 671994
rect 58922 671758 59104 671994
rect 58504 635994 59104 671758
rect 58504 635758 58686 635994
rect 58922 635758 59104 635994
rect 58504 599994 59104 635758
rect 58504 599758 58686 599994
rect 58922 599758 59104 599994
rect 58504 563994 59104 599758
rect 58504 563758 58686 563994
rect 58922 563758 59104 563994
rect 58504 527994 59104 563758
rect 58504 527758 58686 527994
rect 58922 527758 59104 527994
rect 58504 491994 59104 527758
rect 58504 491758 58686 491994
rect 58922 491758 59104 491994
rect 58504 455994 59104 491758
rect 58504 455758 58686 455994
rect 58922 455758 59104 455994
rect 58504 425308 59104 455758
rect 62204 675694 62804 709082
rect 62204 675458 62386 675694
rect 62622 675458 62804 675694
rect 62204 639694 62804 675458
rect 62204 639458 62386 639694
rect 62622 639458 62804 639694
rect 62204 603694 62804 639458
rect 62204 603458 62386 603694
rect 62622 603458 62804 603694
rect 62204 567694 62804 603458
rect 62204 567458 62386 567694
rect 62622 567458 62804 567694
rect 62204 531694 62804 567458
rect 62204 531458 62386 531694
rect 62622 531458 62804 531694
rect 62204 495694 62804 531458
rect 62204 495458 62386 495694
rect 62622 495458 62804 495694
rect 62204 459694 62804 495458
rect 62204 459458 62386 459694
rect 62622 459458 62804 459694
rect 62204 425308 62804 459458
rect 65904 679394 66504 711002
rect 83904 710598 84504 711590
rect 83904 710362 84086 710598
rect 84322 710362 84504 710598
rect 83904 710278 84504 710362
rect 83904 710042 84086 710278
rect 84322 710042 84504 710278
rect 80204 708678 80804 709670
rect 80204 708442 80386 708678
rect 80622 708442 80804 708678
rect 80204 708358 80804 708442
rect 80204 708122 80386 708358
rect 80622 708122 80804 708358
rect 76504 706758 77104 707750
rect 76504 706522 76686 706758
rect 76922 706522 77104 706758
rect 76504 706438 77104 706522
rect 76504 706202 76686 706438
rect 76922 706202 77104 706438
rect 65904 679158 66086 679394
rect 66322 679158 66504 679394
rect 65904 643394 66504 679158
rect 65904 643158 66086 643394
rect 66322 643158 66504 643394
rect 65904 607394 66504 643158
rect 65904 607158 66086 607394
rect 66322 607158 66504 607394
rect 65904 571394 66504 607158
rect 65904 571158 66086 571394
rect 66322 571158 66504 571394
rect 65904 535394 66504 571158
rect 65904 535158 66086 535394
rect 66322 535158 66504 535394
rect 65904 499394 66504 535158
rect 65904 499158 66086 499394
rect 66322 499158 66504 499394
rect 65904 463394 66504 499158
rect 65904 463158 66086 463394
rect 66322 463158 66504 463394
rect 65904 427394 66504 463158
rect 65904 427158 66086 427394
rect 66322 427158 66504 427394
rect 65904 425308 66504 427158
rect 72804 704838 73404 705830
rect 72804 704602 72986 704838
rect 73222 704602 73404 704838
rect 72804 704518 73404 704602
rect 72804 704282 72986 704518
rect 73222 704282 73404 704518
rect 72804 686294 73404 704282
rect 72804 686058 72986 686294
rect 73222 686058 73404 686294
rect 72804 650294 73404 686058
rect 72804 650058 72986 650294
rect 73222 650058 73404 650294
rect 72804 614294 73404 650058
rect 72804 614058 72986 614294
rect 73222 614058 73404 614294
rect 72804 578294 73404 614058
rect 72804 578058 72986 578294
rect 73222 578058 73404 578294
rect 72804 542294 73404 578058
rect 72804 542058 72986 542294
rect 73222 542058 73404 542294
rect 72804 506294 73404 542058
rect 72804 506058 72986 506294
rect 73222 506058 73404 506294
rect 72804 470294 73404 506058
rect 72804 470058 72986 470294
rect 73222 470058 73404 470294
rect 72804 434294 73404 470058
rect 72804 434058 72986 434294
rect 73222 434058 73404 434294
rect 72804 425308 73404 434058
rect 76504 689994 77104 706202
rect 76504 689758 76686 689994
rect 76922 689758 77104 689994
rect 76504 653994 77104 689758
rect 76504 653758 76686 653994
rect 76922 653758 77104 653994
rect 76504 617994 77104 653758
rect 76504 617758 76686 617994
rect 76922 617758 77104 617994
rect 76504 581994 77104 617758
rect 76504 581758 76686 581994
rect 76922 581758 77104 581994
rect 76504 545994 77104 581758
rect 76504 545758 76686 545994
rect 76922 545758 77104 545994
rect 76504 509994 77104 545758
rect 76504 509758 76686 509994
rect 76922 509758 77104 509994
rect 76504 473994 77104 509758
rect 76504 473758 76686 473994
rect 76922 473758 77104 473994
rect 76504 437994 77104 473758
rect 76504 437758 76686 437994
rect 76922 437758 77104 437994
rect 76504 425308 77104 437758
rect 80204 693694 80804 708122
rect 80204 693458 80386 693694
rect 80622 693458 80804 693694
rect 80204 657694 80804 693458
rect 80204 657458 80386 657694
rect 80622 657458 80804 657694
rect 80204 621694 80804 657458
rect 80204 621458 80386 621694
rect 80622 621458 80804 621694
rect 80204 585694 80804 621458
rect 80204 585458 80386 585694
rect 80622 585458 80804 585694
rect 80204 549694 80804 585458
rect 80204 549458 80386 549694
rect 80622 549458 80804 549694
rect 80204 513694 80804 549458
rect 80204 513458 80386 513694
rect 80622 513458 80804 513694
rect 80204 477694 80804 513458
rect 80204 477458 80386 477694
rect 80622 477458 80804 477694
rect 80204 441694 80804 477458
rect 80204 441458 80386 441694
rect 80622 441458 80804 441694
rect 80204 425308 80804 441458
rect 83904 697394 84504 710042
rect 101904 711558 102504 711590
rect 101904 711322 102086 711558
rect 102322 711322 102504 711558
rect 101904 711238 102504 711322
rect 101904 711002 102086 711238
rect 102322 711002 102504 711238
rect 98204 709638 98804 709670
rect 98204 709402 98386 709638
rect 98622 709402 98804 709638
rect 98204 709318 98804 709402
rect 98204 709082 98386 709318
rect 98622 709082 98804 709318
rect 94504 707718 95104 707750
rect 94504 707482 94686 707718
rect 94922 707482 95104 707718
rect 94504 707398 95104 707482
rect 94504 707162 94686 707398
rect 94922 707162 95104 707398
rect 83904 697158 84086 697394
rect 84322 697158 84504 697394
rect 83904 661394 84504 697158
rect 83904 661158 84086 661394
rect 84322 661158 84504 661394
rect 83904 625394 84504 661158
rect 83904 625158 84086 625394
rect 84322 625158 84504 625394
rect 83904 589394 84504 625158
rect 83904 589158 84086 589394
rect 84322 589158 84504 589394
rect 83904 553394 84504 589158
rect 83904 553158 84086 553394
rect 84322 553158 84504 553394
rect 83904 517394 84504 553158
rect 83904 517158 84086 517394
rect 84322 517158 84504 517394
rect 83904 481394 84504 517158
rect 83904 481158 84086 481394
rect 84322 481158 84504 481394
rect 83904 445394 84504 481158
rect 83904 445158 84086 445394
rect 84322 445158 84504 445394
rect 83904 425308 84504 445158
rect 90804 705798 91404 705830
rect 90804 705562 90986 705798
rect 91222 705562 91404 705798
rect 90804 705478 91404 705562
rect 90804 705242 90986 705478
rect 91222 705242 91404 705478
rect 90804 668294 91404 705242
rect 90804 668058 90986 668294
rect 91222 668058 91404 668294
rect 90804 632294 91404 668058
rect 90804 632058 90986 632294
rect 91222 632058 91404 632294
rect 90804 596294 91404 632058
rect 90804 596058 90986 596294
rect 91222 596058 91404 596294
rect 90804 560294 91404 596058
rect 90804 560058 90986 560294
rect 91222 560058 91404 560294
rect 90804 524294 91404 560058
rect 90804 524058 90986 524294
rect 91222 524058 91404 524294
rect 90804 488294 91404 524058
rect 90804 488058 90986 488294
rect 91222 488058 91404 488294
rect 90804 452294 91404 488058
rect 90804 452058 90986 452294
rect 91222 452058 91404 452294
rect 90804 425308 91404 452058
rect 94504 671994 95104 707162
rect 94504 671758 94686 671994
rect 94922 671758 95104 671994
rect 94504 635994 95104 671758
rect 94504 635758 94686 635994
rect 94922 635758 95104 635994
rect 94504 599994 95104 635758
rect 94504 599758 94686 599994
rect 94922 599758 95104 599994
rect 94504 563994 95104 599758
rect 94504 563758 94686 563994
rect 94922 563758 95104 563994
rect 94504 527994 95104 563758
rect 94504 527758 94686 527994
rect 94922 527758 95104 527994
rect 94504 491994 95104 527758
rect 94504 491758 94686 491994
rect 94922 491758 95104 491994
rect 94504 455994 95104 491758
rect 94504 455758 94686 455994
rect 94922 455758 95104 455994
rect 94504 425308 95104 455758
rect 98204 675694 98804 709082
rect 98204 675458 98386 675694
rect 98622 675458 98804 675694
rect 98204 639694 98804 675458
rect 98204 639458 98386 639694
rect 98622 639458 98804 639694
rect 98204 603694 98804 639458
rect 98204 603458 98386 603694
rect 98622 603458 98804 603694
rect 98204 567694 98804 603458
rect 98204 567458 98386 567694
rect 98622 567458 98804 567694
rect 98204 531694 98804 567458
rect 98204 531458 98386 531694
rect 98622 531458 98804 531694
rect 98204 495694 98804 531458
rect 98204 495458 98386 495694
rect 98622 495458 98804 495694
rect 98204 459694 98804 495458
rect 98204 459458 98386 459694
rect 98622 459458 98804 459694
rect 98204 425308 98804 459458
rect 101904 679394 102504 711002
rect 119904 710598 120504 711590
rect 119904 710362 120086 710598
rect 120322 710362 120504 710598
rect 119904 710278 120504 710362
rect 119904 710042 120086 710278
rect 120322 710042 120504 710278
rect 116204 708678 116804 709670
rect 116204 708442 116386 708678
rect 116622 708442 116804 708678
rect 116204 708358 116804 708442
rect 116204 708122 116386 708358
rect 116622 708122 116804 708358
rect 112504 706758 113104 707750
rect 112504 706522 112686 706758
rect 112922 706522 113104 706758
rect 112504 706438 113104 706522
rect 112504 706202 112686 706438
rect 112922 706202 113104 706438
rect 101904 679158 102086 679394
rect 102322 679158 102504 679394
rect 101904 643394 102504 679158
rect 101904 643158 102086 643394
rect 102322 643158 102504 643394
rect 101904 607394 102504 643158
rect 101904 607158 102086 607394
rect 102322 607158 102504 607394
rect 101904 571394 102504 607158
rect 101904 571158 102086 571394
rect 102322 571158 102504 571394
rect 101904 535394 102504 571158
rect 101904 535158 102086 535394
rect 102322 535158 102504 535394
rect 101904 499394 102504 535158
rect 101904 499158 102086 499394
rect 102322 499158 102504 499394
rect 101904 463394 102504 499158
rect 101904 463158 102086 463394
rect 102322 463158 102504 463394
rect 101904 427394 102504 463158
rect 101904 427158 102086 427394
rect 102322 427158 102504 427394
rect 101904 425308 102504 427158
rect 108804 704838 109404 705830
rect 108804 704602 108986 704838
rect 109222 704602 109404 704838
rect 108804 704518 109404 704602
rect 108804 704282 108986 704518
rect 109222 704282 109404 704518
rect 108804 686294 109404 704282
rect 108804 686058 108986 686294
rect 109222 686058 109404 686294
rect 108804 650294 109404 686058
rect 108804 650058 108986 650294
rect 109222 650058 109404 650294
rect 108804 614294 109404 650058
rect 108804 614058 108986 614294
rect 109222 614058 109404 614294
rect 108804 578294 109404 614058
rect 108804 578058 108986 578294
rect 109222 578058 109404 578294
rect 108804 542294 109404 578058
rect 108804 542058 108986 542294
rect 109222 542058 109404 542294
rect 108804 506294 109404 542058
rect 108804 506058 108986 506294
rect 109222 506058 109404 506294
rect 108804 470294 109404 506058
rect 108804 470058 108986 470294
rect 109222 470058 109404 470294
rect 108804 434294 109404 470058
rect 108804 434058 108986 434294
rect 109222 434058 109404 434294
rect 108804 425308 109404 434058
rect 112504 689994 113104 706202
rect 112504 689758 112686 689994
rect 112922 689758 113104 689994
rect 112504 653994 113104 689758
rect 112504 653758 112686 653994
rect 112922 653758 113104 653994
rect 112504 617994 113104 653758
rect 112504 617758 112686 617994
rect 112922 617758 113104 617994
rect 112504 581994 113104 617758
rect 112504 581758 112686 581994
rect 112922 581758 113104 581994
rect 112504 545994 113104 581758
rect 112504 545758 112686 545994
rect 112922 545758 113104 545994
rect 112504 509994 113104 545758
rect 112504 509758 112686 509994
rect 112922 509758 113104 509994
rect 112504 473994 113104 509758
rect 112504 473758 112686 473994
rect 112922 473758 113104 473994
rect 112504 437994 113104 473758
rect 112504 437758 112686 437994
rect 112922 437758 113104 437994
rect 112504 425308 113104 437758
rect 116204 693694 116804 708122
rect 116204 693458 116386 693694
rect 116622 693458 116804 693694
rect 116204 657694 116804 693458
rect 116204 657458 116386 657694
rect 116622 657458 116804 657694
rect 116204 621694 116804 657458
rect 116204 621458 116386 621694
rect 116622 621458 116804 621694
rect 116204 585694 116804 621458
rect 116204 585458 116386 585694
rect 116622 585458 116804 585694
rect 116204 549694 116804 585458
rect 116204 549458 116386 549694
rect 116622 549458 116804 549694
rect 116204 513694 116804 549458
rect 116204 513458 116386 513694
rect 116622 513458 116804 513694
rect 116204 477694 116804 513458
rect 116204 477458 116386 477694
rect 116622 477458 116804 477694
rect 116204 441694 116804 477458
rect 116204 441458 116386 441694
rect 116622 441458 116804 441694
rect 116204 425308 116804 441458
rect 119904 697394 120504 710042
rect 137904 711558 138504 711590
rect 137904 711322 138086 711558
rect 138322 711322 138504 711558
rect 137904 711238 138504 711322
rect 137904 711002 138086 711238
rect 138322 711002 138504 711238
rect 134204 709638 134804 709670
rect 134204 709402 134386 709638
rect 134622 709402 134804 709638
rect 134204 709318 134804 709402
rect 134204 709082 134386 709318
rect 134622 709082 134804 709318
rect 130504 707718 131104 707750
rect 130504 707482 130686 707718
rect 130922 707482 131104 707718
rect 130504 707398 131104 707482
rect 130504 707162 130686 707398
rect 130922 707162 131104 707398
rect 119904 697158 120086 697394
rect 120322 697158 120504 697394
rect 119904 661394 120504 697158
rect 119904 661158 120086 661394
rect 120322 661158 120504 661394
rect 119904 625394 120504 661158
rect 119904 625158 120086 625394
rect 120322 625158 120504 625394
rect 119904 589394 120504 625158
rect 119904 589158 120086 589394
rect 120322 589158 120504 589394
rect 119904 553394 120504 589158
rect 119904 553158 120086 553394
rect 120322 553158 120504 553394
rect 119904 517394 120504 553158
rect 119904 517158 120086 517394
rect 120322 517158 120504 517394
rect 119904 481394 120504 517158
rect 119904 481158 120086 481394
rect 120322 481158 120504 481394
rect 119904 445394 120504 481158
rect 119904 445158 120086 445394
rect 120322 445158 120504 445394
rect 119904 425308 120504 445158
rect 126804 705798 127404 705830
rect 126804 705562 126986 705798
rect 127222 705562 127404 705798
rect 126804 705478 127404 705562
rect 126804 705242 126986 705478
rect 127222 705242 127404 705478
rect 126804 668294 127404 705242
rect 126804 668058 126986 668294
rect 127222 668058 127404 668294
rect 126804 632294 127404 668058
rect 126804 632058 126986 632294
rect 127222 632058 127404 632294
rect 126804 596294 127404 632058
rect 126804 596058 126986 596294
rect 127222 596058 127404 596294
rect 126804 560294 127404 596058
rect 126804 560058 126986 560294
rect 127222 560058 127404 560294
rect 126804 524294 127404 560058
rect 126804 524058 126986 524294
rect 127222 524058 127404 524294
rect 126804 488294 127404 524058
rect 126804 488058 126986 488294
rect 127222 488058 127404 488294
rect 126804 452294 127404 488058
rect 126804 452058 126986 452294
rect 127222 452058 127404 452294
rect 126804 425308 127404 452058
rect 130504 671994 131104 707162
rect 130504 671758 130686 671994
rect 130922 671758 131104 671994
rect 130504 635994 131104 671758
rect 130504 635758 130686 635994
rect 130922 635758 131104 635994
rect 130504 599994 131104 635758
rect 130504 599758 130686 599994
rect 130922 599758 131104 599994
rect 130504 563994 131104 599758
rect 130504 563758 130686 563994
rect 130922 563758 131104 563994
rect 130504 527994 131104 563758
rect 130504 527758 130686 527994
rect 130922 527758 131104 527994
rect 130504 491994 131104 527758
rect 130504 491758 130686 491994
rect 130922 491758 131104 491994
rect 130504 455994 131104 491758
rect 130504 455758 130686 455994
rect 130922 455758 131104 455994
rect 130504 425308 131104 455758
rect 134204 675694 134804 709082
rect 134204 675458 134386 675694
rect 134622 675458 134804 675694
rect 134204 639694 134804 675458
rect 134204 639458 134386 639694
rect 134622 639458 134804 639694
rect 134204 603694 134804 639458
rect 134204 603458 134386 603694
rect 134622 603458 134804 603694
rect 134204 567694 134804 603458
rect 134204 567458 134386 567694
rect 134622 567458 134804 567694
rect 134204 531694 134804 567458
rect 134204 531458 134386 531694
rect 134622 531458 134804 531694
rect 134204 495694 134804 531458
rect 134204 495458 134386 495694
rect 134622 495458 134804 495694
rect 134204 459694 134804 495458
rect 134204 459458 134386 459694
rect 134622 459458 134804 459694
rect 134204 425308 134804 459458
rect 137904 679394 138504 711002
rect 155904 710598 156504 711590
rect 155904 710362 156086 710598
rect 156322 710362 156504 710598
rect 155904 710278 156504 710362
rect 155904 710042 156086 710278
rect 156322 710042 156504 710278
rect 152204 708678 152804 709670
rect 152204 708442 152386 708678
rect 152622 708442 152804 708678
rect 152204 708358 152804 708442
rect 152204 708122 152386 708358
rect 152622 708122 152804 708358
rect 148504 706758 149104 707750
rect 148504 706522 148686 706758
rect 148922 706522 149104 706758
rect 148504 706438 149104 706522
rect 148504 706202 148686 706438
rect 148922 706202 149104 706438
rect 137904 679158 138086 679394
rect 138322 679158 138504 679394
rect 137904 643394 138504 679158
rect 137904 643158 138086 643394
rect 138322 643158 138504 643394
rect 137904 607394 138504 643158
rect 137904 607158 138086 607394
rect 138322 607158 138504 607394
rect 137904 571394 138504 607158
rect 137904 571158 138086 571394
rect 138322 571158 138504 571394
rect 137904 535394 138504 571158
rect 137904 535158 138086 535394
rect 138322 535158 138504 535394
rect 137904 499394 138504 535158
rect 137904 499158 138086 499394
rect 138322 499158 138504 499394
rect 137904 463394 138504 499158
rect 137904 463158 138086 463394
rect 138322 463158 138504 463394
rect 137904 427394 138504 463158
rect 137904 427158 138086 427394
rect 138322 427158 138504 427394
rect 137904 425308 138504 427158
rect 144804 704838 145404 705830
rect 144804 704602 144986 704838
rect 145222 704602 145404 704838
rect 144804 704518 145404 704602
rect 144804 704282 144986 704518
rect 145222 704282 145404 704518
rect 144804 686294 145404 704282
rect 144804 686058 144986 686294
rect 145222 686058 145404 686294
rect 144804 650294 145404 686058
rect 144804 650058 144986 650294
rect 145222 650058 145404 650294
rect 144804 614294 145404 650058
rect 144804 614058 144986 614294
rect 145222 614058 145404 614294
rect 144804 578294 145404 614058
rect 144804 578058 144986 578294
rect 145222 578058 145404 578294
rect 144804 542294 145404 578058
rect 144804 542058 144986 542294
rect 145222 542058 145404 542294
rect 144804 506294 145404 542058
rect 144804 506058 144986 506294
rect 145222 506058 145404 506294
rect 144804 470294 145404 506058
rect 144804 470058 144986 470294
rect 145222 470058 145404 470294
rect 144804 434294 145404 470058
rect 144804 434058 144986 434294
rect 145222 434058 145404 434294
rect 144804 425308 145404 434058
rect 148504 689994 149104 706202
rect 148504 689758 148686 689994
rect 148922 689758 149104 689994
rect 148504 653994 149104 689758
rect 148504 653758 148686 653994
rect 148922 653758 149104 653994
rect 148504 617994 149104 653758
rect 148504 617758 148686 617994
rect 148922 617758 149104 617994
rect 148504 581994 149104 617758
rect 148504 581758 148686 581994
rect 148922 581758 149104 581994
rect 148504 545994 149104 581758
rect 148504 545758 148686 545994
rect 148922 545758 149104 545994
rect 148504 509994 149104 545758
rect 148504 509758 148686 509994
rect 148922 509758 149104 509994
rect 148504 473994 149104 509758
rect 148504 473758 148686 473994
rect 148922 473758 149104 473994
rect 148504 437994 149104 473758
rect 148504 437758 148686 437994
rect 148922 437758 149104 437994
rect 148504 425308 149104 437758
rect 152204 693694 152804 708122
rect 152204 693458 152386 693694
rect 152622 693458 152804 693694
rect 152204 657694 152804 693458
rect 152204 657458 152386 657694
rect 152622 657458 152804 657694
rect 152204 621694 152804 657458
rect 152204 621458 152386 621694
rect 152622 621458 152804 621694
rect 152204 585694 152804 621458
rect 152204 585458 152386 585694
rect 152622 585458 152804 585694
rect 152204 549694 152804 585458
rect 152204 549458 152386 549694
rect 152622 549458 152804 549694
rect 152204 513694 152804 549458
rect 152204 513458 152386 513694
rect 152622 513458 152804 513694
rect 152204 477694 152804 513458
rect 152204 477458 152386 477694
rect 152622 477458 152804 477694
rect 152204 441694 152804 477458
rect 152204 441458 152386 441694
rect 152622 441458 152804 441694
rect 152204 425308 152804 441458
rect 155904 697394 156504 710042
rect 173904 711558 174504 711590
rect 173904 711322 174086 711558
rect 174322 711322 174504 711558
rect 173904 711238 174504 711322
rect 173904 711002 174086 711238
rect 174322 711002 174504 711238
rect 170204 709638 170804 709670
rect 170204 709402 170386 709638
rect 170622 709402 170804 709638
rect 170204 709318 170804 709402
rect 170204 709082 170386 709318
rect 170622 709082 170804 709318
rect 166504 707718 167104 707750
rect 166504 707482 166686 707718
rect 166922 707482 167104 707718
rect 166504 707398 167104 707482
rect 166504 707162 166686 707398
rect 166922 707162 167104 707398
rect 155904 697158 156086 697394
rect 156322 697158 156504 697394
rect 155904 661394 156504 697158
rect 155904 661158 156086 661394
rect 156322 661158 156504 661394
rect 155904 625394 156504 661158
rect 155904 625158 156086 625394
rect 156322 625158 156504 625394
rect 155904 589394 156504 625158
rect 155904 589158 156086 589394
rect 156322 589158 156504 589394
rect 155904 553394 156504 589158
rect 155904 553158 156086 553394
rect 156322 553158 156504 553394
rect 155904 517394 156504 553158
rect 155904 517158 156086 517394
rect 156322 517158 156504 517394
rect 155904 481394 156504 517158
rect 155904 481158 156086 481394
rect 156322 481158 156504 481394
rect 155904 445394 156504 481158
rect 155904 445158 156086 445394
rect 156322 445158 156504 445394
rect 155904 425308 156504 445158
rect 162804 705798 163404 705830
rect 162804 705562 162986 705798
rect 163222 705562 163404 705798
rect 162804 705478 163404 705562
rect 162804 705242 162986 705478
rect 163222 705242 163404 705478
rect 162804 668294 163404 705242
rect 162804 668058 162986 668294
rect 163222 668058 163404 668294
rect 162804 632294 163404 668058
rect 162804 632058 162986 632294
rect 163222 632058 163404 632294
rect 162804 596294 163404 632058
rect 162804 596058 162986 596294
rect 163222 596058 163404 596294
rect 162804 560294 163404 596058
rect 162804 560058 162986 560294
rect 163222 560058 163404 560294
rect 162804 524294 163404 560058
rect 162804 524058 162986 524294
rect 163222 524058 163404 524294
rect 162804 488294 163404 524058
rect 162804 488058 162986 488294
rect 163222 488058 163404 488294
rect 162804 452294 163404 488058
rect 162804 452058 162986 452294
rect 163222 452058 163404 452294
rect 162804 425308 163404 452058
rect 166504 671994 167104 707162
rect 166504 671758 166686 671994
rect 166922 671758 167104 671994
rect 166504 635994 167104 671758
rect 166504 635758 166686 635994
rect 166922 635758 167104 635994
rect 166504 599994 167104 635758
rect 166504 599758 166686 599994
rect 166922 599758 167104 599994
rect 166504 563994 167104 599758
rect 166504 563758 166686 563994
rect 166922 563758 167104 563994
rect 166504 527994 167104 563758
rect 166504 527758 166686 527994
rect 166922 527758 167104 527994
rect 166504 491994 167104 527758
rect 166504 491758 166686 491994
rect 166922 491758 167104 491994
rect 166504 455994 167104 491758
rect 166504 455758 166686 455994
rect 166922 455758 167104 455994
rect 166504 425308 167104 455758
rect 170204 675694 170804 709082
rect 170204 675458 170386 675694
rect 170622 675458 170804 675694
rect 170204 639694 170804 675458
rect 170204 639458 170386 639694
rect 170622 639458 170804 639694
rect 170204 603694 170804 639458
rect 170204 603458 170386 603694
rect 170622 603458 170804 603694
rect 170204 567694 170804 603458
rect 170204 567458 170386 567694
rect 170622 567458 170804 567694
rect 170204 531694 170804 567458
rect 170204 531458 170386 531694
rect 170622 531458 170804 531694
rect 170204 495694 170804 531458
rect 170204 495458 170386 495694
rect 170622 495458 170804 495694
rect 170204 459694 170804 495458
rect 170204 459458 170386 459694
rect 170622 459458 170804 459694
rect 170204 425308 170804 459458
rect 173904 679394 174504 711002
rect 191904 710598 192504 711590
rect 191904 710362 192086 710598
rect 192322 710362 192504 710598
rect 191904 710278 192504 710362
rect 191904 710042 192086 710278
rect 192322 710042 192504 710278
rect 188204 708678 188804 709670
rect 188204 708442 188386 708678
rect 188622 708442 188804 708678
rect 188204 708358 188804 708442
rect 188204 708122 188386 708358
rect 188622 708122 188804 708358
rect 184504 706758 185104 707750
rect 184504 706522 184686 706758
rect 184922 706522 185104 706758
rect 184504 706438 185104 706522
rect 184504 706202 184686 706438
rect 184922 706202 185104 706438
rect 173904 679158 174086 679394
rect 174322 679158 174504 679394
rect 173904 643394 174504 679158
rect 173904 643158 174086 643394
rect 174322 643158 174504 643394
rect 173904 607394 174504 643158
rect 173904 607158 174086 607394
rect 174322 607158 174504 607394
rect 173904 571394 174504 607158
rect 173904 571158 174086 571394
rect 174322 571158 174504 571394
rect 173904 535394 174504 571158
rect 173904 535158 174086 535394
rect 174322 535158 174504 535394
rect 173904 499394 174504 535158
rect 173904 499158 174086 499394
rect 174322 499158 174504 499394
rect 173904 463394 174504 499158
rect 173904 463158 174086 463394
rect 174322 463158 174504 463394
rect 173904 427394 174504 463158
rect 173904 427158 174086 427394
rect 174322 427158 174504 427394
rect 173904 425308 174504 427158
rect 180804 704838 181404 705830
rect 180804 704602 180986 704838
rect 181222 704602 181404 704838
rect 180804 704518 181404 704602
rect 180804 704282 180986 704518
rect 181222 704282 181404 704518
rect 180804 686294 181404 704282
rect 180804 686058 180986 686294
rect 181222 686058 181404 686294
rect 180804 650294 181404 686058
rect 180804 650058 180986 650294
rect 181222 650058 181404 650294
rect 180804 614294 181404 650058
rect 180804 614058 180986 614294
rect 181222 614058 181404 614294
rect 180804 578294 181404 614058
rect 180804 578058 180986 578294
rect 181222 578058 181404 578294
rect 180804 542294 181404 578058
rect 180804 542058 180986 542294
rect 181222 542058 181404 542294
rect 180804 506294 181404 542058
rect 180804 506058 180986 506294
rect 181222 506058 181404 506294
rect 180804 470294 181404 506058
rect 180804 470058 180986 470294
rect 181222 470058 181404 470294
rect 180804 434294 181404 470058
rect 180804 434058 180986 434294
rect 181222 434058 181404 434294
rect 40272 416294 40620 416476
rect 40272 416058 40328 416294
rect 40564 416058 40620 416294
rect 40272 415876 40620 416058
rect 176000 416294 176348 416476
rect 176000 416058 176056 416294
rect 176292 416058 176348 416294
rect 176000 415876 176348 416058
rect 36804 398058 36986 398294
rect 37222 398058 37404 398294
rect 36804 362294 37404 398058
rect 40952 398294 41300 398476
rect 40952 398058 41008 398294
rect 41244 398058 41300 398294
rect 40952 397876 41300 398058
rect 175320 398294 175668 398476
rect 175320 398058 175376 398294
rect 175612 398058 175668 398294
rect 175320 397876 175668 398058
rect 180804 398294 181404 434058
rect 180804 398058 180986 398294
rect 181222 398058 181404 398294
rect 40272 380294 40620 380476
rect 40272 380058 40328 380294
rect 40564 380058 40620 380294
rect 40272 379876 40620 380058
rect 176000 380294 176348 380476
rect 176000 380058 176056 380294
rect 176292 380058 176348 380294
rect 176000 379876 176348 380058
rect 36804 362058 36986 362294
rect 37222 362058 37404 362294
rect 36804 326294 37404 362058
rect 40952 362294 41300 362476
rect 40952 362058 41008 362294
rect 41244 362058 41300 362294
rect 40952 361876 41300 362058
rect 175320 362294 175668 362476
rect 175320 362058 175376 362294
rect 175612 362058 175668 362294
rect 175320 361876 175668 362058
rect 180804 362294 181404 398058
rect 180804 362058 180986 362294
rect 181222 362058 181404 362294
rect 40272 344294 40620 344476
rect 40272 344058 40328 344294
rect 40564 344058 40620 344294
rect 40272 343876 40620 344058
rect 176000 344294 176348 344476
rect 176000 344058 176056 344294
rect 176292 344058 176348 344294
rect 176000 343876 176348 344058
rect 93534 340076 93622 340136
rect 56056 339690 56116 340000
rect 57144 339690 57204 340000
rect 58232 339690 58292 340000
rect 59592 339690 59652 340000
rect 55998 339630 56116 339690
rect 57102 339630 57204 339690
rect 58206 339630 58292 339690
rect 59494 339630 59652 339690
rect 60544 339690 60604 340000
rect 61768 339690 61828 340000
rect 63128 339690 63188 340000
rect 64216 339690 64276 340000
rect 65440 339690 65500 340000
rect 60544 339630 60658 339690
rect 61768 339630 61946 339690
rect 63128 339630 63234 339690
rect 64216 339630 64338 339690
rect 36804 326058 36986 326294
rect 37222 326058 37404 326294
rect 36804 290294 37404 326058
rect 36804 290058 36986 290294
rect 37222 290058 37404 290294
rect 36804 254294 37404 290058
rect 36804 254058 36986 254294
rect 37222 254058 37404 254294
rect 36804 218294 37404 254058
rect 40504 329994 41104 338000
rect 40504 329758 40686 329994
rect 40922 329758 41104 329994
rect 40504 293994 41104 329758
rect 40504 293758 40686 293994
rect 40922 293758 41104 293994
rect 40504 257994 41104 293758
rect 40504 257758 40686 257994
rect 40922 257758 41104 257994
rect 40504 243568 41104 257758
rect 44204 333694 44804 338000
rect 47715 337788 47781 337789
rect 47715 337724 47716 337788
rect 47780 337724 47781 337788
rect 47715 337723 47781 337724
rect 44204 333458 44386 333694
rect 44622 333458 44804 333694
rect 44204 297694 44804 333458
rect 44204 297458 44386 297694
rect 44622 297458 44804 297694
rect 44204 261694 44804 297458
rect 44204 261458 44386 261694
rect 44622 261458 44804 261694
rect 44204 243568 44804 261458
rect 42563 242996 42629 242997
rect 42563 242932 42564 242996
rect 42628 242932 42629 242996
rect 42563 242931 42629 242932
rect 36804 218058 36986 218294
rect 37222 218058 37404 218294
rect 36804 182294 37404 218058
rect 36804 182058 36986 182294
rect 37222 182058 37404 182294
rect 36804 146294 37404 182058
rect 36804 146058 36986 146294
rect 37222 146058 37404 146294
rect 36804 110294 37404 146058
rect 36804 110058 36986 110294
rect 37222 110058 37404 110294
rect 36804 74294 37404 110058
rect 36804 74058 36986 74294
rect 37222 74058 37404 74294
rect 36804 38294 37404 74058
rect 42566 39949 42626 242931
rect 44208 218294 44528 218476
rect 44208 218058 44250 218294
rect 44486 218058 44528 218294
rect 44208 217876 44528 218058
rect 44208 182294 44528 182476
rect 44208 182058 44250 182294
rect 44486 182058 44528 182294
rect 44208 181876 44528 182058
rect 44208 146294 44528 146476
rect 44208 146058 44250 146294
rect 44486 146058 44528 146294
rect 44208 145876 44528 146058
rect 44208 110294 44528 110476
rect 44208 110058 44250 110294
rect 44486 110058 44528 110294
rect 44208 109876 44528 110058
rect 44208 74294 44528 74476
rect 44208 74058 44250 74294
rect 44486 74058 44528 74294
rect 44208 73876 44528 74058
rect 42563 39948 42629 39949
rect 42563 39884 42564 39948
rect 42628 39884 42629 39948
rect 42563 39883 42629 39884
rect 47718 38589 47778 337723
rect 47904 337394 48504 338000
rect 47904 337158 48086 337394
rect 48322 337158 48504 337394
rect 47904 301394 48504 337158
rect 47904 301158 48086 301394
rect 48322 301158 48504 301394
rect 47904 265394 48504 301158
rect 47904 265158 48086 265394
rect 48322 265158 48504 265394
rect 47904 243568 48504 265158
rect 54804 308294 55404 338000
rect 55998 337925 56058 339630
rect 55995 337924 56061 337925
rect 55995 337860 55996 337924
rect 56060 337860 56061 337924
rect 55995 337859 56061 337860
rect 57102 337517 57162 339630
rect 58206 337653 58266 339630
rect 58203 337652 58269 337653
rect 58203 337588 58204 337652
rect 58268 337588 58269 337652
rect 58203 337587 58269 337588
rect 57099 337516 57165 337517
rect 57099 337452 57100 337516
rect 57164 337452 57165 337516
rect 57099 337451 57165 337452
rect 54804 308058 54986 308294
rect 55222 308058 55404 308294
rect 54804 272294 55404 308058
rect 54804 272058 54986 272294
rect 55222 272058 55404 272294
rect 54804 243568 55404 272058
rect 58504 311994 59104 338000
rect 59494 337245 59554 339630
rect 60598 337381 60658 339630
rect 61886 337653 61946 339630
rect 61883 337652 61949 337653
rect 61883 337588 61884 337652
rect 61948 337588 61949 337652
rect 61883 337587 61949 337588
rect 60595 337380 60661 337381
rect 60595 337316 60596 337380
rect 60660 337316 60661 337380
rect 60595 337315 60661 337316
rect 59491 337244 59557 337245
rect 59491 337180 59492 337244
rect 59556 337180 59557 337244
rect 59491 337179 59557 337180
rect 58504 311758 58686 311994
rect 58922 311758 59104 311994
rect 58504 275994 59104 311758
rect 58504 275758 58686 275994
rect 58922 275758 59104 275994
rect 58504 243568 59104 275758
rect 62204 315694 62804 338000
rect 63174 337653 63234 339630
rect 63171 337652 63237 337653
rect 63171 337588 63172 337652
rect 63236 337588 63237 337652
rect 63171 337587 63237 337588
rect 64278 337517 64338 339630
rect 65382 339630 65500 339690
rect 66528 339690 66588 340000
rect 67616 339690 67676 340000
rect 66528 339630 66730 339690
rect 65382 337653 65442 339630
rect 65379 337652 65445 337653
rect 65379 337588 65380 337652
rect 65444 337588 65445 337652
rect 65379 337587 65445 337588
rect 64275 337516 64341 337517
rect 64275 337452 64276 337516
rect 64340 337452 64341 337516
rect 64275 337451 64341 337452
rect 62204 315458 62386 315694
rect 62622 315458 62804 315694
rect 62204 279694 62804 315458
rect 62204 279458 62386 279694
rect 62622 279458 62804 279694
rect 62204 243568 62804 279458
rect 65904 319394 66504 338000
rect 66670 337653 66730 339630
rect 67590 339630 67676 339690
rect 68296 339690 68356 340000
rect 68704 339690 68764 340000
rect 70064 339690 70124 340000
rect 70744 339690 70804 340000
rect 71288 339690 71348 340000
rect 72376 339690 72436 340000
rect 68296 339630 68386 339690
rect 67590 337789 67650 339630
rect 68326 337925 68386 339630
rect 68694 339630 68764 339690
rect 69982 339630 70124 339690
rect 70718 339630 70804 339690
rect 71270 339630 71348 339690
rect 72374 339630 72436 339690
rect 73464 339690 73524 340000
rect 73600 339690 73660 340000
rect 74552 339690 74612 340000
rect 75912 339690 75972 340000
rect 73464 339630 73538 339690
rect 73600 339630 73722 339690
rect 74552 339630 74642 339690
rect 68323 337924 68389 337925
rect 68323 337860 68324 337924
rect 68388 337860 68389 337924
rect 68323 337859 68389 337860
rect 67587 337788 67653 337789
rect 67587 337724 67588 337788
rect 67652 337724 67653 337788
rect 67587 337723 67653 337724
rect 68694 337653 68754 339630
rect 66667 337652 66733 337653
rect 66667 337588 66668 337652
rect 66732 337588 66733 337652
rect 66667 337587 66733 337588
rect 68691 337652 68757 337653
rect 68691 337588 68692 337652
rect 68756 337588 68757 337652
rect 68691 337587 68757 337588
rect 69982 337381 70042 339630
rect 70718 337653 70778 339630
rect 71270 337789 71330 339630
rect 71267 337788 71333 337789
rect 71267 337724 71268 337788
rect 71332 337724 71333 337788
rect 71267 337723 71333 337724
rect 70715 337652 70781 337653
rect 70715 337588 70716 337652
rect 70780 337588 70781 337652
rect 70715 337587 70781 337588
rect 72374 337517 72434 339630
rect 72371 337516 72437 337517
rect 72371 337452 72372 337516
rect 72436 337452 72437 337516
rect 72371 337451 72437 337452
rect 69979 337380 70045 337381
rect 69979 337316 69980 337380
rect 70044 337316 70045 337380
rect 69979 337315 70045 337316
rect 65904 319158 66086 319394
rect 66322 319158 66504 319394
rect 65904 283394 66504 319158
rect 65904 283158 66086 283394
rect 66322 283158 66504 283394
rect 65904 247394 66504 283158
rect 65904 247158 66086 247394
rect 66322 247158 66504 247394
rect 65904 243568 66504 247158
rect 72804 326294 73404 338000
rect 73478 337789 73538 339630
rect 73475 337788 73541 337789
rect 73475 337724 73476 337788
rect 73540 337724 73541 337788
rect 73475 337723 73541 337724
rect 73662 337653 73722 339630
rect 74582 337653 74642 339630
rect 75870 339630 75972 339690
rect 76048 339690 76108 340000
rect 77000 339690 77060 340000
rect 78088 339690 78148 340000
rect 78496 339690 78556 340000
rect 76048 339630 76114 339690
rect 75870 337789 75930 339630
rect 75867 337788 75933 337789
rect 75867 337724 75868 337788
rect 75932 337724 75933 337788
rect 75867 337723 75933 337724
rect 73659 337652 73725 337653
rect 73659 337588 73660 337652
rect 73724 337588 73725 337652
rect 73659 337587 73725 337588
rect 74579 337652 74645 337653
rect 74579 337588 74580 337652
rect 74644 337588 74645 337652
rect 74579 337587 74645 337588
rect 76054 336837 76114 339630
rect 76974 339630 77060 339690
rect 78078 339630 78148 339690
rect 78446 339630 78556 339690
rect 79448 339690 79508 340000
rect 80672 339690 80732 340000
rect 81080 339690 81140 340000
rect 81760 339690 81820 340000
rect 79448 339630 79610 339690
rect 80672 339630 80898 339690
rect 81080 339630 81266 339690
rect 76974 338197 77034 339630
rect 76971 338196 77037 338197
rect 76971 338132 76972 338196
rect 77036 338132 77037 338196
rect 76971 338131 77037 338132
rect 76051 336836 76117 336837
rect 76051 336772 76052 336836
rect 76116 336772 76117 336836
rect 76051 336771 76117 336772
rect 72804 326058 72986 326294
rect 73222 326058 73404 326294
rect 72804 290294 73404 326058
rect 72804 290058 72986 290294
rect 73222 290058 73404 290294
rect 72804 254294 73404 290058
rect 72804 254058 72986 254294
rect 73222 254058 73404 254294
rect 72804 243568 73404 254058
rect 76504 329994 77104 338000
rect 78078 337925 78138 339630
rect 78075 337924 78141 337925
rect 78075 337860 78076 337924
rect 78140 337860 78141 337924
rect 78075 337859 78141 337860
rect 78446 337653 78506 339630
rect 79550 337653 79610 339630
rect 80838 338330 80898 339630
rect 80838 338270 81082 338330
rect 78443 337652 78509 337653
rect 78443 337588 78444 337652
rect 78508 337588 78509 337652
rect 78443 337587 78509 337588
rect 79547 337652 79613 337653
rect 79547 337588 79548 337652
rect 79612 337588 79613 337652
rect 79547 337587 79613 337588
rect 76504 329758 76686 329994
rect 76922 329758 77104 329994
rect 76504 293994 77104 329758
rect 76504 293758 76686 293994
rect 76922 293758 77104 293994
rect 76504 257994 77104 293758
rect 76504 257758 76686 257994
rect 76922 257758 77104 257994
rect 76504 243568 77104 257758
rect 80204 333694 80804 338000
rect 81022 337653 81082 338270
rect 81019 337652 81085 337653
rect 81019 337588 81020 337652
rect 81084 337588 81085 337652
rect 81019 337587 81085 337588
rect 81206 336837 81266 339630
rect 81758 339630 81820 339690
rect 82848 339690 82908 340000
rect 83528 339690 83588 340000
rect 83936 339690 83996 340000
rect 85296 339690 85356 340000
rect 82848 339630 82922 339690
rect 81758 337653 81818 339630
rect 82862 337789 82922 339630
rect 83414 339630 83588 339690
rect 83782 339630 83996 339690
rect 85254 339630 85356 339690
rect 85976 339690 86036 340000
rect 86384 339690 86444 340000
rect 85976 339630 86050 339690
rect 82859 337788 82925 337789
rect 82859 337724 82860 337788
rect 82924 337724 82925 337788
rect 82859 337723 82925 337724
rect 83414 337653 83474 339630
rect 81755 337652 81821 337653
rect 81755 337588 81756 337652
rect 81820 337588 81821 337652
rect 81755 337587 81821 337588
rect 83411 337652 83477 337653
rect 83411 337588 83412 337652
rect 83476 337588 83477 337652
rect 83411 337587 83477 337588
rect 83595 336972 83661 336973
rect 83595 336908 83596 336972
rect 83660 336970 83661 336972
rect 83782 336970 83842 339630
rect 83660 336910 83842 336970
rect 83904 337394 84504 338000
rect 85254 337653 85314 339630
rect 85251 337652 85317 337653
rect 85251 337588 85252 337652
rect 85316 337588 85317 337652
rect 85251 337587 85317 337588
rect 83904 337158 84086 337394
rect 84322 337158 84504 337394
rect 85990 337381 86050 339630
rect 86358 339630 86444 339690
rect 87608 339690 87668 340000
rect 88288 339690 88348 340000
rect 87608 339630 87706 339690
rect 86358 337653 86418 339630
rect 87646 337789 87706 339630
rect 88198 339630 88348 339690
rect 88696 339690 88756 340000
rect 89784 339690 89844 340000
rect 91008 339690 91068 340000
rect 88696 339630 88810 339690
rect 89784 339630 89914 339690
rect 87643 337788 87709 337789
rect 87643 337724 87644 337788
rect 87708 337724 87709 337788
rect 87643 337723 87709 337724
rect 88198 337653 88258 339630
rect 88750 337653 88810 339630
rect 89854 337653 89914 339630
rect 90958 339630 91068 339690
rect 91144 339690 91204 340000
rect 92232 339690 92292 340000
rect 93320 339690 93380 340000
rect 91144 339630 91570 339690
rect 92232 339630 92306 339690
rect 93320 339630 93410 339690
rect 90958 338197 91018 339630
rect 90955 338196 91021 338197
rect 90955 338132 90956 338196
rect 91020 338132 91021 338196
rect 90955 338131 91021 338132
rect 86355 337652 86421 337653
rect 86355 337588 86356 337652
rect 86420 337588 86421 337652
rect 86355 337587 86421 337588
rect 88195 337652 88261 337653
rect 88195 337588 88196 337652
rect 88260 337588 88261 337652
rect 88195 337587 88261 337588
rect 88747 337652 88813 337653
rect 88747 337588 88748 337652
rect 88812 337588 88813 337652
rect 88747 337587 88813 337588
rect 89851 337652 89917 337653
rect 89851 337588 89852 337652
rect 89916 337588 89917 337652
rect 89851 337587 89917 337588
rect 85987 337380 86053 337381
rect 85987 337316 85988 337380
rect 86052 337316 86053 337380
rect 85987 337315 86053 337316
rect 83660 336908 83661 336910
rect 83595 336907 83661 336908
rect 81203 336836 81269 336837
rect 81203 336772 81204 336836
rect 81268 336772 81269 336836
rect 81203 336771 81269 336772
rect 80204 333458 80386 333694
rect 80622 333458 80804 333694
rect 80204 297694 80804 333458
rect 80204 297458 80386 297694
rect 80622 297458 80804 297694
rect 80204 261694 80804 297458
rect 80204 261458 80386 261694
rect 80622 261458 80804 261694
rect 80204 243568 80804 261458
rect 83904 301394 84504 337158
rect 83904 301158 84086 301394
rect 84322 301158 84504 301394
rect 83904 265394 84504 301158
rect 83904 265158 84086 265394
rect 84322 265158 84504 265394
rect 83904 243568 84504 265158
rect 90804 308294 91404 338000
rect 91510 337789 91570 339630
rect 91507 337788 91573 337789
rect 91507 337724 91508 337788
rect 91572 337724 91573 337788
rect 91507 337723 91573 337724
rect 92246 337653 92306 339630
rect 93350 337789 93410 339630
rect 93347 337788 93413 337789
rect 93347 337724 93348 337788
rect 93412 337724 93413 337788
rect 93347 337723 93413 337724
rect 93534 337653 93594 340076
rect 94408 339690 94468 340000
rect 95768 339690 95828 340000
rect 94270 339630 94468 339690
rect 95742 339630 95828 339690
rect 96040 339690 96100 340000
rect 96992 339690 97052 340000
rect 98080 339690 98140 340000
rect 96040 339630 96170 339690
rect 96992 339630 97090 339690
rect 94270 337789 94330 339630
rect 94267 337788 94333 337789
rect 94267 337724 94268 337788
rect 94332 337724 94333 337788
rect 94267 337723 94333 337724
rect 92243 337652 92309 337653
rect 92243 337588 92244 337652
rect 92308 337588 92309 337652
rect 92243 337587 92309 337588
rect 93531 337652 93597 337653
rect 93531 337588 93532 337652
rect 93596 337588 93597 337652
rect 93531 337587 93597 337588
rect 90804 308058 90986 308294
rect 91222 308058 91404 308294
rect 90804 272294 91404 308058
rect 90804 272058 90986 272294
rect 91222 272058 91404 272294
rect 90804 243568 91404 272058
rect 94504 311994 95104 338000
rect 95742 337653 95802 339630
rect 95739 337652 95805 337653
rect 95739 337588 95740 337652
rect 95804 337588 95805 337652
rect 95739 337587 95805 337588
rect 96110 336837 96170 339630
rect 97030 337653 97090 339630
rect 97950 339630 98140 339690
rect 98488 339690 98548 340000
rect 99168 339690 99228 340000
rect 100936 339690 100996 340000
rect 103520 339690 103580 340000
rect 98488 339630 98930 339690
rect 97950 337925 98010 339630
rect 97947 337924 98013 337925
rect 97947 337860 97948 337924
rect 98012 337860 98013 337924
rect 97947 337859 98013 337860
rect 97027 337652 97093 337653
rect 97027 337588 97028 337652
rect 97092 337588 97093 337652
rect 97027 337587 97093 337588
rect 96107 336836 96173 336837
rect 96107 336772 96108 336836
rect 96172 336772 96173 336836
rect 96107 336771 96173 336772
rect 94504 311758 94686 311994
rect 94922 311758 95104 311994
rect 94504 275994 95104 311758
rect 94504 275758 94686 275994
rect 94922 275758 95104 275994
rect 94504 243568 95104 275758
rect 98204 315694 98804 338000
rect 98870 336837 98930 339630
rect 99054 339630 99228 339690
rect 100894 339630 100996 339690
rect 103286 339630 103580 339690
rect 105968 339690 106028 340000
rect 108280 339690 108340 340000
rect 105968 339630 106106 339690
rect 99054 337789 99114 339630
rect 99051 337788 99117 337789
rect 99051 337724 99052 337788
rect 99116 337724 99117 337788
rect 99051 337723 99117 337724
rect 100894 337653 100954 339630
rect 100891 337652 100957 337653
rect 100891 337588 100892 337652
rect 100956 337588 100957 337652
rect 100891 337587 100957 337588
rect 98867 336836 98933 336837
rect 98867 336772 98868 336836
rect 98932 336772 98933 336836
rect 98867 336771 98933 336772
rect 98204 315458 98386 315694
rect 98622 315458 98804 315694
rect 98204 279694 98804 315458
rect 98204 279458 98386 279694
rect 98622 279458 98804 279694
rect 98204 243568 98804 279458
rect 101904 319394 102504 338000
rect 103286 336834 103346 339630
rect 106046 337653 106106 339630
rect 108254 339630 108340 339690
rect 111000 339690 111060 340000
rect 113448 339690 113508 340000
rect 111000 339630 111074 339690
rect 108254 337653 108314 339630
rect 106043 337652 106109 337653
rect 106043 337588 106044 337652
rect 106108 337588 106109 337652
rect 106043 337587 106109 337588
rect 108251 337652 108317 337653
rect 108251 337588 108252 337652
rect 108316 337588 108317 337652
rect 108251 337587 108317 337588
rect 103467 336836 103533 336837
rect 103467 336834 103468 336836
rect 103286 336774 103468 336834
rect 103467 336772 103468 336774
rect 103532 336772 103533 336836
rect 103467 336771 103533 336772
rect 101904 319158 102086 319394
rect 102322 319158 102504 319394
rect 101904 283394 102504 319158
rect 101904 283158 102086 283394
rect 102322 283158 102504 283394
rect 101904 247394 102504 283158
rect 101904 247158 102086 247394
rect 102322 247158 102504 247394
rect 101904 243568 102504 247158
rect 108804 326294 109404 338000
rect 111014 337653 111074 339630
rect 113406 339630 113508 339690
rect 115896 339690 115956 340000
rect 118480 339690 118540 340000
rect 120928 339690 120988 340000
rect 123512 339690 123572 340000
rect 125960 339690 126020 340000
rect 128544 339690 128604 340000
rect 115896 339630 116042 339690
rect 118480 339630 118618 339690
rect 120928 339630 121010 339690
rect 123512 339630 123586 339690
rect 111011 337652 111077 337653
rect 111011 337588 111012 337652
rect 111076 337588 111077 337652
rect 111011 337587 111077 337588
rect 108804 326058 108986 326294
rect 109222 326058 109404 326294
rect 108804 290294 109404 326058
rect 108804 290058 108986 290294
rect 109222 290058 109404 290294
rect 108804 254294 109404 290058
rect 108804 254058 108986 254294
rect 109222 254058 109404 254294
rect 108804 243568 109404 254058
rect 112504 329994 113104 338000
rect 113406 337653 113466 339630
rect 113403 337652 113469 337653
rect 113403 337588 113404 337652
rect 113468 337588 113469 337652
rect 113403 337587 113469 337588
rect 115982 337245 116042 339630
rect 115979 337244 116045 337245
rect 115979 337180 115980 337244
rect 116044 337180 116045 337244
rect 115979 337179 116045 337180
rect 112504 329758 112686 329994
rect 112922 329758 113104 329994
rect 112504 293994 113104 329758
rect 112504 293758 112686 293994
rect 112922 293758 113104 293994
rect 112504 257994 113104 293758
rect 112504 257758 112686 257994
rect 112922 257758 113104 257994
rect 112504 243568 113104 257758
rect 116204 333694 116804 338000
rect 118558 337653 118618 339630
rect 118555 337652 118621 337653
rect 118555 337588 118556 337652
rect 118620 337588 118621 337652
rect 118555 337587 118621 337588
rect 116204 333458 116386 333694
rect 116622 333458 116804 333694
rect 116204 297694 116804 333458
rect 116204 297458 116386 297694
rect 116622 297458 116804 297694
rect 116204 261694 116804 297458
rect 116204 261458 116386 261694
rect 116622 261458 116804 261694
rect 116204 243568 116804 261458
rect 119904 337394 120504 338000
rect 120950 337653 121010 339630
rect 123526 337653 123586 339630
rect 125918 339630 126020 339690
rect 128494 339630 128604 339690
rect 130992 339690 131052 340000
rect 133440 339690 133500 340000
rect 135888 339690 135948 340000
rect 130992 339630 131130 339690
rect 133440 339630 133522 339690
rect 125918 337653 125978 339630
rect 120947 337652 121013 337653
rect 120947 337588 120948 337652
rect 121012 337588 121013 337652
rect 120947 337587 121013 337588
rect 123523 337652 123589 337653
rect 123523 337588 123524 337652
rect 123588 337588 123589 337652
rect 123523 337587 123589 337588
rect 125915 337652 125981 337653
rect 125915 337588 125916 337652
rect 125980 337588 125981 337652
rect 125915 337587 125981 337588
rect 119904 337158 120086 337394
rect 120322 337158 120504 337394
rect 119904 301394 120504 337158
rect 119904 301158 120086 301394
rect 120322 301158 120504 301394
rect 119904 265394 120504 301158
rect 119904 265158 120086 265394
rect 120322 265158 120504 265394
rect 119904 243568 120504 265158
rect 126804 308294 127404 338000
rect 128494 337653 128554 339630
rect 131070 338197 131130 339630
rect 131067 338196 131133 338197
rect 131067 338132 131068 338196
rect 131132 338132 131133 338196
rect 131067 338131 131133 338132
rect 128491 337652 128557 337653
rect 128491 337588 128492 337652
rect 128556 337588 128557 337652
rect 128491 337587 128557 337588
rect 126804 308058 126986 308294
rect 127222 308058 127404 308294
rect 126804 272294 127404 308058
rect 126804 272058 126986 272294
rect 127222 272058 127404 272294
rect 126804 243568 127404 272058
rect 130504 311994 131104 338000
rect 133462 337653 133522 339630
rect 135854 339630 135948 339690
rect 138472 339690 138532 340000
rect 140920 339690 140980 340000
rect 143368 339690 143428 340000
rect 145952 339690 146012 340000
rect 138472 339630 138674 339690
rect 140920 339630 141066 339690
rect 143368 339630 143458 339690
rect 145952 339630 146034 339690
rect 133459 337652 133525 337653
rect 133459 337588 133460 337652
rect 133524 337588 133525 337652
rect 133459 337587 133525 337588
rect 130504 311758 130686 311994
rect 130922 311758 131104 311994
rect 130504 275994 131104 311758
rect 130504 275758 130686 275994
rect 130922 275758 131104 275994
rect 130504 243568 131104 275758
rect 134204 315694 134804 338000
rect 135854 337653 135914 339630
rect 135851 337652 135917 337653
rect 135851 337588 135852 337652
rect 135916 337588 135917 337652
rect 135851 337587 135917 337588
rect 134204 315458 134386 315694
rect 134622 315458 134804 315694
rect 134204 279694 134804 315458
rect 134204 279458 134386 279694
rect 134622 279458 134804 279694
rect 134204 243568 134804 279458
rect 137904 319394 138504 338000
rect 138614 337653 138674 339630
rect 141006 337653 141066 339630
rect 143398 337789 143458 339630
rect 143395 337788 143461 337789
rect 143395 337724 143396 337788
rect 143460 337724 143461 337788
rect 143395 337723 143461 337724
rect 138611 337652 138677 337653
rect 138611 337588 138612 337652
rect 138676 337588 138677 337652
rect 138611 337587 138677 337588
rect 141003 337652 141069 337653
rect 141003 337588 141004 337652
rect 141068 337588 141069 337652
rect 141003 337587 141069 337588
rect 137904 319158 138086 319394
rect 138322 319158 138504 319394
rect 137904 283394 138504 319158
rect 137904 283158 138086 283394
rect 138322 283158 138504 283394
rect 137904 247394 138504 283158
rect 137904 247158 138086 247394
rect 138322 247158 138504 247394
rect 137904 243568 138504 247158
rect 144804 326294 145404 338000
rect 145974 337653 146034 339630
rect 145971 337652 146037 337653
rect 145971 337588 145972 337652
rect 146036 337588 146037 337652
rect 145971 337587 146037 337588
rect 144804 326058 144986 326294
rect 145222 326058 145404 326294
rect 144804 290294 145404 326058
rect 144804 290058 144986 290294
rect 145222 290058 145404 290294
rect 144804 254294 145404 290058
rect 144804 254058 144986 254294
rect 145222 254058 145404 254294
rect 144804 243568 145404 254058
rect 148504 329994 149104 338000
rect 148504 329758 148686 329994
rect 148922 329758 149104 329994
rect 148504 293994 149104 329758
rect 148504 293758 148686 293994
rect 148922 293758 149104 293994
rect 148504 257994 149104 293758
rect 148504 257758 148686 257994
rect 148922 257758 149104 257994
rect 148504 243568 149104 257758
rect 152204 333694 152804 338000
rect 152204 333458 152386 333694
rect 152622 333458 152804 333694
rect 152204 297694 152804 333458
rect 152204 297458 152386 297694
rect 152622 297458 152804 297694
rect 152204 261694 152804 297458
rect 152204 261458 152386 261694
rect 152622 261458 152804 261694
rect 152204 243568 152804 261458
rect 155904 337394 156504 338000
rect 155904 337158 156086 337394
rect 156322 337158 156504 337394
rect 155904 301394 156504 337158
rect 155904 301158 156086 301394
rect 156322 301158 156504 301394
rect 155904 265394 156504 301158
rect 155904 265158 156086 265394
rect 156322 265158 156504 265394
rect 155904 243568 156504 265158
rect 162804 308294 163404 338000
rect 162804 308058 162986 308294
rect 163222 308058 163404 308294
rect 162804 272294 163404 308058
rect 162804 272058 162986 272294
rect 163222 272058 163404 272294
rect 162804 243568 163404 272058
rect 166504 311994 167104 338000
rect 166504 311758 166686 311994
rect 166922 311758 167104 311994
rect 166504 275994 167104 311758
rect 166504 275758 166686 275994
rect 166922 275758 167104 275994
rect 166504 243568 167104 275758
rect 170204 315694 170804 338000
rect 170204 315458 170386 315694
rect 170622 315458 170804 315694
rect 170204 279694 170804 315458
rect 170204 279458 170386 279694
rect 170622 279458 170804 279694
rect 170204 243568 170804 279458
rect 173904 319394 174504 338000
rect 173904 319158 174086 319394
rect 174322 319158 174504 319394
rect 173904 283394 174504 319158
rect 173904 283158 174086 283394
rect 174322 283158 174504 283394
rect 173904 247394 174504 283158
rect 173904 247158 174086 247394
rect 174322 247158 174504 247394
rect 173904 243568 174504 247158
rect 180804 326294 181404 362058
rect 180804 326058 180986 326294
rect 181222 326058 181404 326294
rect 180804 290294 181404 326058
rect 180804 290058 180986 290294
rect 181222 290058 181404 290294
rect 180804 254294 181404 290058
rect 180804 254058 180986 254294
rect 181222 254058 181404 254294
rect 180804 243568 181404 254058
rect 184504 689994 185104 706202
rect 184504 689758 184686 689994
rect 184922 689758 185104 689994
rect 184504 653994 185104 689758
rect 184504 653758 184686 653994
rect 184922 653758 185104 653994
rect 184504 617994 185104 653758
rect 184504 617758 184686 617994
rect 184922 617758 185104 617994
rect 184504 581994 185104 617758
rect 184504 581758 184686 581994
rect 184922 581758 185104 581994
rect 184504 545994 185104 581758
rect 184504 545758 184686 545994
rect 184922 545758 185104 545994
rect 184504 509994 185104 545758
rect 184504 509758 184686 509994
rect 184922 509758 185104 509994
rect 184504 473994 185104 509758
rect 184504 473758 184686 473994
rect 184922 473758 185104 473994
rect 184504 437994 185104 473758
rect 184504 437758 184686 437994
rect 184922 437758 185104 437994
rect 184504 401994 185104 437758
rect 184504 401758 184686 401994
rect 184922 401758 185104 401994
rect 184504 365994 185104 401758
rect 184504 365758 184686 365994
rect 184922 365758 185104 365994
rect 184504 329994 185104 365758
rect 184504 329758 184686 329994
rect 184922 329758 185104 329994
rect 184504 293994 185104 329758
rect 184504 293758 184686 293994
rect 184922 293758 185104 293994
rect 184504 257994 185104 293758
rect 184504 257758 184686 257994
rect 184922 257758 185104 257994
rect 184504 243568 185104 257758
rect 188204 693694 188804 708122
rect 188204 693458 188386 693694
rect 188622 693458 188804 693694
rect 188204 657694 188804 693458
rect 188204 657458 188386 657694
rect 188622 657458 188804 657694
rect 188204 621694 188804 657458
rect 188204 621458 188386 621694
rect 188622 621458 188804 621694
rect 188204 585694 188804 621458
rect 188204 585458 188386 585694
rect 188622 585458 188804 585694
rect 188204 549694 188804 585458
rect 188204 549458 188386 549694
rect 188622 549458 188804 549694
rect 188204 513694 188804 549458
rect 188204 513458 188386 513694
rect 188622 513458 188804 513694
rect 188204 477694 188804 513458
rect 188204 477458 188386 477694
rect 188622 477458 188804 477694
rect 188204 441694 188804 477458
rect 188204 441458 188386 441694
rect 188622 441458 188804 441694
rect 188204 405694 188804 441458
rect 188204 405458 188386 405694
rect 188622 405458 188804 405694
rect 188204 369694 188804 405458
rect 188204 369458 188386 369694
rect 188622 369458 188804 369694
rect 188204 333694 188804 369458
rect 188204 333458 188386 333694
rect 188622 333458 188804 333694
rect 188204 297694 188804 333458
rect 188204 297458 188386 297694
rect 188622 297458 188804 297694
rect 188204 261694 188804 297458
rect 188204 261458 188386 261694
rect 188622 261458 188804 261694
rect 188204 243568 188804 261458
rect 191904 697394 192504 710042
rect 209904 711558 210504 711590
rect 209904 711322 210086 711558
rect 210322 711322 210504 711558
rect 209904 711238 210504 711322
rect 209904 711002 210086 711238
rect 210322 711002 210504 711238
rect 206204 709638 206804 709670
rect 206204 709402 206386 709638
rect 206622 709402 206804 709638
rect 206204 709318 206804 709402
rect 206204 709082 206386 709318
rect 206622 709082 206804 709318
rect 202504 707718 203104 707750
rect 202504 707482 202686 707718
rect 202922 707482 203104 707718
rect 202504 707398 203104 707482
rect 202504 707162 202686 707398
rect 202922 707162 203104 707398
rect 191904 697158 192086 697394
rect 192322 697158 192504 697394
rect 191904 661394 192504 697158
rect 191904 661158 192086 661394
rect 192322 661158 192504 661394
rect 191904 625394 192504 661158
rect 191904 625158 192086 625394
rect 192322 625158 192504 625394
rect 191904 589394 192504 625158
rect 191904 589158 192086 589394
rect 192322 589158 192504 589394
rect 191904 553394 192504 589158
rect 191904 553158 192086 553394
rect 192322 553158 192504 553394
rect 191904 517394 192504 553158
rect 191904 517158 192086 517394
rect 192322 517158 192504 517394
rect 191904 481394 192504 517158
rect 191904 481158 192086 481394
rect 192322 481158 192504 481394
rect 191904 445394 192504 481158
rect 191904 445158 192086 445394
rect 192322 445158 192504 445394
rect 191904 409394 192504 445158
rect 191904 409158 192086 409394
rect 192322 409158 192504 409394
rect 191904 373394 192504 409158
rect 191904 373158 192086 373394
rect 192322 373158 192504 373394
rect 191904 337394 192504 373158
rect 191904 337158 192086 337394
rect 192322 337158 192504 337394
rect 191904 301394 192504 337158
rect 191904 301158 192086 301394
rect 192322 301158 192504 301394
rect 191904 265394 192504 301158
rect 191904 265158 192086 265394
rect 192322 265158 192504 265394
rect 191904 243568 192504 265158
rect 198804 705798 199404 705830
rect 198804 705562 198986 705798
rect 199222 705562 199404 705798
rect 198804 705478 199404 705562
rect 198804 705242 198986 705478
rect 199222 705242 199404 705478
rect 198804 668294 199404 705242
rect 198804 668058 198986 668294
rect 199222 668058 199404 668294
rect 198804 632294 199404 668058
rect 198804 632058 198986 632294
rect 199222 632058 199404 632294
rect 198804 596294 199404 632058
rect 198804 596058 198986 596294
rect 199222 596058 199404 596294
rect 198804 560294 199404 596058
rect 198804 560058 198986 560294
rect 199222 560058 199404 560294
rect 198804 524294 199404 560058
rect 198804 524058 198986 524294
rect 199222 524058 199404 524294
rect 198804 488294 199404 524058
rect 198804 488058 198986 488294
rect 199222 488058 199404 488294
rect 198804 452294 199404 488058
rect 198804 452058 198986 452294
rect 199222 452058 199404 452294
rect 198804 416294 199404 452058
rect 198804 416058 198986 416294
rect 199222 416058 199404 416294
rect 198804 380294 199404 416058
rect 198804 380058 198986 380294
rect 199222 380058 199404 380294
rect 198804 344294 199404 380058
rect 198804 344058 198986 344294
rect 199222 344058 199404 344294
rect 198804 308294 199404 344058
rect 198804 308058 198986 308294
rect 199222 308058 199404 308294
rect 198804 272294 199404 308058
rect 198804 272058 198986 272294
rect 199222 272058 199404 272294
rect 198804 243568 199404 272058
rect 202504 671994 203104 707162
rect 202504 671758 202686 671994
rect 202922 671758 203104 671994
rect 202504 635994 203104 671758
rect 202504 635758 202686 635994
rect 202922 635758 203104 635994
rect 202504 599994 203104 635758
rect 202504 599758 202686 599994
rect 202922 599758 203104 599994
rect 202504 563994 203104 599758
rect 202504 563758 202686 563994
rect 202922 563758 203104 563994
rect 202504 527994 203104 563758
rect 202504 527758 202686 527994
rect 202922 527758 203104 527994
rect 202504 491994 203104 527758
rect 202504 491758 202686 491994
rect 202922 491758 203104 491994
rect 202504 455994 203104 491758
rect 202504 455758 202686 455994
rect 202922 455758 203104 455994
rect 202504 419994 203104 455758
rect 202504 419758 202686 419994
rect 202922 419758 203104 419994
rect 202504 383994 203104 419758
rect 202504 383758 202686 383994
rect 202922 383758 203104 383994
rect 202504 347994 203104 383758
rect 202504 347758 202686 347994
rect 202922 347758 203104 347994
rect 202504 311994 203104 347758
rect 202504 311758 202686 311994
rect 202922 311758 203104 311994
rect 202504 275994 203104 311758
rect 202504 275758 202686 275994
rect 202922 275758 203104 275994
rect 202504 243568 203104 275758
rect 206204 675694 206804 709082
rect 206204 675458 206386 675694
rect 206622 675458 206804 675694
rect 206204 639694 206804 675458
rect 206204 639458 206386 639694
rect 206622 639458 206804 639694
rect 206204 603694 206804 639458
rect 206204 603458 206386 603694
rect 206622 603458 206804 603694
rect 206204 567694 206804 603458
rect 206204 567458 206386 567694
rect 206622 567458 206804 567694
rect 206204 531694 206804 567458
rect 206204 531458 206386 531694
rect 206622 531458 206804 531694
rect 206204 495694 206804 531458
rect 206204 495458 206386 495694
rect 206622 495458 206804 495694
rect 206204 459694 206804 495458
rect 206204 459458 206386 459694
rect 206622 459458 206804 459694
rect 206204 423694 206804 459458
rect 206204 423458 206386 423694
rect 206622 423458 206804 423694
rect 206204 387694 206804 423458
rect 206204 387458 206386 387694
rect 206622 387458 206804 387694
rect 206204 351694 206804 387458
rect 206204 351458 206386 351694
rect 206622 351458 206804 351694
rect 206204 315694 206804 351458
rect 206204 315458 206386 315694
rect 206622 315458 206804 315694
rect 206204 279694 206804 315458
rect 206204 279458 206386 279694
rect 206622 279458 206804 279694
rect 206204 243568 206804 279458
rect 209904 679394 210504 711002
rect 227904 710598 228504 711590
rect 227904 710362 228086 710598
rect 228322 710362 228504 710598
rect 227904 710278 228504 710362
rect 227904 710042 228086 710278
rect 228322 710042 228504 710278
rect 224204 708678 224804 709670
rect 224204 708442 224386 708678
rect 224622 708442 224804 708678
rect 224204 708358 224804 708442
rect 224204 708122 224386 708358
rect 224622 708122 224804 708358
rect 220504 706758 221104 707750
rect 220504 706522 220686 706758
rect 220922 706522 221104 706758
rect 220504 706438 221104 706522
rect 220504 706202 220686 706438
rect 220922 706202 221104 706438
rect 209904 679158 210086 679394
rect 210322 679158 210504 679394
rect 209904 643394 210504 679158
rect 209904 643158 210086 643394
rect 210322 643158 210504 643394
rect 209904 607394 210504 643158
rect 209904 607158 210086 607394
rect 210322 607158 210504 607394
rect 209904 571394 210504 607158
rect 209904 571158 210086 571394
rect 210322 571158 210504 571394
rect 209904 535394 210504 571158
rect 209904 535158 210086 535394
rect 210322 535158 210504 535394
rect 209904 499394 210504 535158
rect 209904 499158 210086 499394
rect 210322 499158 210504 499394
rect 209904 463394 210504 499158
rect 209904 463158 210086 463394
rect 210322 463158 210504 463394
rect 209904 427394 210504 463158
rect 209904 427158 210086 427394
rect 210322 427158 210504 427394
rect 209904 391394 210504 427158
rect 209904 391158 210086 391394
rect 210322 391158 210504 391394
rect 209904 355394 210504 391158
rect 209904 355158 210086 355394
rect 210322 355158 210504 355394
rect 209904 319394 210504 355158
rect 209904 319158 210086 319394
rect 210322 319158 210504 319394
rect 209904 283394 210504 319158
rect 209904 283158 210086 283394
rect 210322 283158 210504 283394
rect 209904 247394 210504 283158
rect 209904 247158 210086 247394
rect 210322 247158 210504 247394
rect 209904 243568 210504 247158
rect 216804 704838 217404 705830
rect 216804 704602 216986 704838
rect 217222 704602 217404 704838
rect 216804 704518 217404 704602
rect 216804 704282 216986 704518
rect 217222 704282 217404 704518
rect 216804 686294 217404 704282
rect 216804 686058 216986 686294
rect 217222 686058 217404 686294
rect 216804 650294 217404 686058
rect 216804 650058 216986 650294
rect 217222 650058 217404 650294
rect 216804 614294 217404 650058
rect 216804 614058 216986 614294
rect 217222 614058 217404 614294
rect 216804 578294 217404 614058
rect 216804 578058 216986 578294
rect 217222 578058 217404 578294
rect 216804 542294 217404 578058
rect 216804 542058 216986 542294
rect 217222 542058 217404 542294
rect 216804 506294 217404 542058
rect 216804 506058 216986 506294
rect 217222 506058 217404 506294
rect 216804 470294 217404 506058
rect 216804 470058 216986 470294
rect 217222 470058 217404 470294
rect 216804 434294 217404 470058
rect 216804 434058 216986 434294
rect 217222 434058 217404 434294
rect 216804 398294 217404 434058
rect 216804 398058 216986 398294
rect 217222 398058 217404 398294
rect 216804 362294 217404 398058
rect 216804 362058 216986 362294
rect 217222 362058 217404 362294
rect 216804 326294 217404 362058
rect 216804 326058 216986 326294
rect 217222 326058 217404 326294
rect 216804 290294 217404 326058
rect 216804 290058 216986 290294
rect 217222 290058 217404 290294
rect 216804 254294 217404 290058
rect 216804 254058 216986 254294
rect 217222 254058 217404 254294
rect 216804 243568 217404 254058
rect 220504 689994 221104 706202
rect 220504 689758 220686 689994
rect 220922 689758 221104 689994
rect 220504 653994 221104 689758
rect 220504 653758 220686 653994
rect 220922 653758 221104 653994
rect 220504 617994 221104 653758
rect 220504 617758 220686 617994
rect 220922 617758 221104 617994
rect 220504 581994 221104 617758
rect 220504 581758 220686 581994
rect 220922 581758 221104 581994
rect 220504 545994 221104 581758
rect 220504 545758 220686 545994
rect 220922 545758 221104 545994
rect 220504 509994 221104 545758
rect 220504 509758 220686 509994
rect 220922 509758 221104 509994
rect 220504 473994 221104 509758
rect 220504 473758 220686 473994
rect 220922 473758 221104 473994
rect 220504 437994 221104 473758
rect 220504 437758 220686 437994
rect 220922 437758 221104 437994
rect 220504 401994 221104 437758
rect 220504 401758 220686 401994
rect 220922 401758 221104 401994
rect 220504 365994 221104 401758
rect 220504 365758 220686 365994
rect 220922 365758 221104 365994
rect 220504 329994 221104 365758
rect 220504 329758 220686 329994
rect 220922 329758 221104 329994
rect 220504 293994 221104 329758
rect 220504 293758 220686 293994
rect 220922 293758 221104 293994
rect 220504 257994 221104 293758
rect 220504 257758 220686 257994
rect 220922 257758 221104 257994
rect 220504 243568 221104 257758
rect 224204 693694 224804 708122
rect 224204 693458 224386 693694
rect 224622 693458 224804 693694
rect 224204 657694 224804 693458
rect 224204 657458 224386 657694
rect 224622 657458 224804 657694
rect 224204 621694 224804 657458
rect 224204 621458 224386 621694
rect 224622 621458 224804 621694
rect 224204 585694 224804 621458
rect 224204 585458 224386 585694
rect 224622 585458 224804 585694
rect 224204 549694 224804 585458
rect 224204 549458 224386 549694
rect 224622 549458 224804 549694
rect 224204 513694 224804 549458
rect 224204 513458 224386 513694
rect 224622 513458 224804 513694
rect 224204 477694 224804 513458
rect 224204 477458 224386 477694
rect 224622 477458 224804 477694
rect 224204 441694 224804 477458
rect 224204 441458 224386 441694
rect 224622 441458 224804 441694
rect 224204 405694 224804 441458
rect 224204 405458 224386 405694
rect 224622 405458 224804 405694
rect 224204 369694 224804 405458
rect 224204 369458 224386 369694
rect 224622 369458 224804 369694
rect 224204 333694 224804 369458
rect 224204 333458 224386 333694
rect 224622 333458 224804 333694
rect 224204 297694 224804 333458
rect 224204 297458 224386 297694
rect 224622 297458 224804 297694
rect 224204 261694 224804 297458
rect 224204 261458 224386 261694
rect 224622 261458 224804 261694
rect 224204 243568 224804 261458
rect 227904 697394 228504 710042
rect 245904 711558 246504 711590
rect 245904 711322 246086 711558
rect 246322 711322 246504 711558
rect 245904 711238 246504 711322
rect 245904 711002 246086 711238
rect 246322 711002 246504 711238
rect 242204 709638 242804 709670
rect 242204 709402 242386 709638
rect 242622 709402 242804 709638
rect 242204 709318 242804 709402
rect 242204 709082 242386 709318
rect 242622 709082 242804 709318
rect 238504 707718 239104 707750
rect 238504 707482 238686 707718
rect 238922 707482 239104 707718
rect 238504 707398 239104 707482
rect 238504 707162 238686 707398
rect 238922 707162 239104 707398
rect 227904 697158 228086 697394
rect 228322 697158 228504 697394
rect 227904 661394 228504 697158
rect 227904 661158 228086 661394
rect 228322 661158 228504 661394
rect 227904 625394 228504 661158
rect 227904 625158 228086 625394
rect 228322 625158 228504 625394
rect 227904 589394 228504 625158
rect 227904 589158 228086 589394
rect 228322 589158 228504 589394
rect 227904 553394 228504 589158
rect 227904 553158 228086 553394
rect 228322 553158 228504 553394
rect 227904 517394 228504 553158
rect 227904 517158 228086 517394
rect 228322 517158 228504 517394
rect 227904 481394 228504 517158
rect 227904 481158 228086 481394
rect 228322 481158 228504 481394
rect 227904 445394 228504 481158
rect 227904 445158 228086 445394
rect 228322 445158 228504 445394
rect 227904 409394 228504 445158
rect 227904 409158 228086 409394
rect 228322 409158 228504 409394
rect 227904 373394 228504 409158
rect 227904 373158 228086 373394
rect 228322 373158 228504 373394
rect 227904 337394 228504 373158
rect 227904 337158 228086 337394
rect 228322 337158 228504 337394
rect 227904 301394 228504 337158
rect 227904 301158 228086 301394
rect 228322 301158 228504 301394
rect 227904 265394 228504 301158
rect 227904 265158 228086 265394
rect 228322 265158 228504 265394
rect 227904 243568 228504 265158
rect 234804 705798 235404 705830
rect 234804 705562 234986 705798
rect 235222 705562 235404 705798
rect 234804 705478 235404 705562
rect 234804 705242 234986 705478
rect 235222 705242 235404 705478
rect 234804 668294 235404 705242
rect 234804 668058 234986 668294
rect 235222 668058 235404 668294
rect 234804 632294 235404 668058
rect 234804 632058 234986 632294
rect 235222 632058 235404 632294
rect 234804 596294 235404 632058
rect 234804 596058 234986 596294
rect 235222 596058 235404 596294
rect 234804 560294 235404 596058
rect 234804 560058 234986 560294
rect 235222 560058 235404 560294
rect 234804 524294 235404 560058
rect 234804 524058 234986 524294
rect 235222 524058 235404 524294
rect 234804 488294 235404 524058
rect 234804 488058 234986 488294
rect 235222 488058 235404 488294
rect 234804 452294 235404 488058
rect 234804 452058 234986 452294
rect 235222 452058 235404 452294
rect 234804 416294 235404 452058
rect 234804 416058 234986 416294
rect 235222 416058 235404 416294
rect 234804 380294 235404 416058
rect 234804 380058 234986 380294
rect 235222 380058 235404 380294
rect 234804 344294 235404 380058
rect 234804 344058 234986 344294
rect 235222 344058 235404 344294
rect 234804 308294 235404 344058
rect 238504 671994 239104 707162
rect 238504 671758 238686 671994
rect 238922 671758 239104 671994
rect 238504 635994 239104 671758
rect 238504 635758 238686 635994
rect 238922 635758 239104 635994
rect 238504 599994 239104 635758
rect 238504 599758 238686 599994
rect 238922 599758 239104 599994
rect 238504 563994 239104 599758
rect 238504 563758 238686 563994
rect 238922 563758 239104 563994
rect 238504 527994 239104 563758
rect 238504 527758 238686 527994
rect 238922 527758 239104 527994
rect 238504 491994 239104 527758
rect 238504 491758 238686 491994
rect 238922 491758 239104 491994
rect 238504 455994 239104 491758
rect 238504 455758 238686 455994
rect 238922 455758 239104 455994
rect 238504 419994 239104 455758
rect 238504 419758 238686 419994
rect 238922 419758 239104 419994
rect 238504 383994 239104 419758
rect 238504 383758 238686 383994
rect 238922 383758 239104 383994
rect 238504 347994 239104 383758
rect 238504 347758 238686 347994
rect 238922 347758 239104 347994
rect 237419 337380 237485 337381
rect 237419 337316 237420 337380
rect 237484 337316 237485 337380
rect 237419 337315 237485 337316
rect 234804 308058 234986 308294
rect 235222 308058 235404 308294
rect 234804 272294 235404 308058
rect 234804 272058 234986 272294
rect 235222 272058 235404 272294
rect 234804 243568 235404 272058
rect 59568 236294 59888 236476
rect 59568 236058 59610 236294
rect 59846 236058 59888 236294
rect 59568 235876 59888 236058
rect 90288 236294 90608 236476
rect 90288 236058 90330 236294
rect 90566 236058 90608 236294
rect 90288 235876 90608 236058
rect 121008 236294 121328 236476
rect 121008 236058 121050 236294
rect 121286 236058 121328 236294
rect 121008 235876 121328 236058
rect 151728 236294 152048 236476
rect 151728 236058 151770 236294
rect 152006 236058 152048 236294
rect 151728 235876 152048 236058
rect 182448 236294 182768 236476
rect 182448 236058 182490 236294
rect 182726 236058 182768 236294
rect 182448 235876 182768 236058
rect 213168 236294 213488 236476
rect 213168 236058 213210 236294
rect 213446 236058 213488 236294
rect 213168 235876 213488 236058
rect 74928 218294 75248 218476
rect 74928 218058 74970 218294
rect 75206 218058 75248 218294
rect 74928 217876 75248 218058
rect 105648 218294 105968 218476
rect 105648 218058 105690 218294
rect 105926 218058 105968 218294
rect 105648 217876 105968 218058
rect 136368 218294 136688 218476
rect 136368 218058 136410 218294
rect 136646 218058 136688 218294
rect 136368 217876 136688 218058
rect 167088 218294 167408 218476
rect 167088 218058 167130 218294
rect 167366 218058 167408 218294
rect 167088 217876 167408 218058
rect 197808 218294 198128 218476
rect 197808 218058 197850 218294
rect 198086 218058 198128 218294
rect 197808 217876 198128 218058
rect 228528 218294 228848 218476
rect 228528 218058 228570 218294
rect 228806 218058 228848 218294
rect 228528 217876 228848 218058
rect 59568 200294 59888 200476
rect 59568 200058 59610 200294
rect 59846 200058 59888 200294
rect 59568 199876 59888 200058
rect 90288 200294 90608 200476
rect 90288 200058 90330 200294
rect 90566 200058 90608 200294
rect 90288 199876 90608 200058
rect 121008 200294 121328 200476
rect 121008 200058 121050 200294
rect 121286 200058 121328 200294
rect 121008 199876 121328 200058
rect 151728 200294 152048 200476
rect 151728 200058 151770 200294
rect 152006 200058 152048 200294
rect 151728 199876 152048 200058
rect 182448 200294 182768 200476
rect 182448 200058 182490 200294
rect 182726 200058 182768 200294
rect 182448 199876 182768 200058
rect 213168 200294 213488 200476
rect 213168 200058 213210 200294
rect 213446 200058 213488 200294
rect 213168 199876 213488 200058
rect 74928 182294 75248 182476
rect 74928 182058 74970 182294
rect 75206 182058 75248 182294
rect 74928 181876 75248 182058
rect 105648 182294 105968 182476
rect 105648 182058 105690 182294
rect 105926 182058 105968 182294
rect 105648 181876 105968 182058
rect 136368 182294 136688 182476
rect 136368 182058 136410 182294
rect 136646 182058 136688 182294
rect 136368 181876 136688 182058
rect 167088 182294 167408 182476
rect 167088 182058 167130 182294
rect 167366 182058 167408 182294
rect 167088 181876 167408 182058
rect 197808 182294 198128 182476
rect 197808 182058 197850 182294
rect 198086 182058 198128 182294
rect 197808 181876 198128 182058
rect 228528 182294 228848 182476
rect 228528 182058 228570 182294
rect 228806 182058 228848 182294
rect 228528 181876 228848 182058
rect 59568 164294 59888 164476
rect 59568 164058 59610 164294
rect 59846 164058 59888 164294
rect 59568 163876 59888 164058
rect 90288 164294 90608 164476
rect 90288 164058 90330 164294
rect 90566 164058 90608 164294
rect 90288 163876 90608 164058
rect 121008 164294 121328 164476
rect 121008 164058 121050 164294
rect 121286 164058 121328 164294
rect 121008 163876 121328 164058
rect 151728 164294 152048 164476
rect 151728 164058 151770 164294
rect 152006 164058 152048 164294
rect 151728 163876 152048 164058
rect 182448 164294 182768 164476
rect 182448 164058 182490 164294
rect 182726 164058 182768 164294
rect 182448 163876 182768 164058
rect 213168 164294 213488 164476
rect 213168 164058 213210 164294
rect 213446 164058 213488 164294
rect 213168 163876 213488 164058
rect 74928 146294 75248 146476
rect 74928 146058 74970 146294
rect 75206 146058 75248 146294
rect 74928 145876 75248 146058
rect 105648 146294 105968 146476
rect 105648 146058 105690 146294
rect 105926 146058 105968 146294
rect 105648 145876 105968 146058
rect 136368 146294 136688 146476
rect 136368 146058 136410 146294
rect 136646 146058 136688 146294
rect 136368 145876 136688 146058
rect 167088 146294 167408 146476
rect 167088 146058 167130 146294
rect 167366 146058 167408 146294
rect 167088 145876 167408 146058
rect 197808 146294 198128 146476
rect 197808 146058 197850 146294
rect 198086 146058 198128 146294
rect 197808 145876 198128 146058
rect 228528 146294 228848 146476
rect 228528 146058 228570 146294
rect 228806 146058 228848 146294
rect 228528 145876 228848 146058
rect 59568 128294 59888 128476
rect 59568 128058 59610 128294
rect 59846 128058 59888 128294
rect 59568 127876 59888 128058
rect 90288 128294 90608 128476
rect 90288 128058 90330 128294
rect 90566 128058 90608 128294
rect 90288 127876 90608 128058
rect 121008 128294 121328 128476
rect 121008 128058 121050 128294
rect 121286 128058 121328 128294
rect 121008 127876 121328 128058
rect 151728 128294 152048 128476
rect 151728 128058 151770 128294
rect 152006 128058 152048 128294
rect 151728 127876 152048 128058
rect 182448 128294 182768 128476
rect 182448 128058 182490 128294
rect 182726 128058 182768 128294
rect 182448 127876 182768 128058
rect 213168 128294 213488 128476
rect 213168 128058 213210 128294
rect 213446 128058 213488 128294
rect 213168 127876 213488 128058
rect 74928 110294 75248 110476
rect 74928 110058 74970 110294
rect 75206 110058 75248 110294
rect 74928 109876 75248 110058
rect 105648 110294 105968 110476
rect 105648 110058 105690 110294
rect 105926 110058 105968 110294
rect 105648 109876 105968 110058
rect 136368 110294 136688 110476
rect 136368 110058 136410 110294
rect 136646 110058 136688 110294
rect 136368 109876 136688 110058
rect 167088 110294 167408 110476
rect 167088 110058 167130 110294
rect 167366 110058 167408 110294
rect 167088 109876 167408 110058
rect 197808 110294 198128 110476
rect 197808 110058 197850 110294
rect 198086 110058 198128 110294
rect 197808 109876 198128 110058
rect 228528 110294 228848 110476
rect 228528 110058 228570 110294
rect 228806 110058 228848 110294
rect 228528 109876 228848 110058
rect 59568 92294 59888 92476
rect 59568 92058 59610 92294
rect 59846 92058 59888 92294
rect 59568 91876 59888 92058
rect 90288 92294 90608 92476
rect 90288 92058 90330 92294
rect 90566 92058 90608 92294
rect 90288 91876 90608 92058
rect 121008 92294 121328 92476
rect 121008 92058 121050 92294
rect 121286 92058 121328 92294
rect 121008 91876 121328 92058
rect 151728 92294 152048 92476
rect 151728 92058 151770 92294
rect 152006 92058 152048 92294
rect 151728 91876 152048 92058
rect 182448 92294 182768 92476
rect 182448 92058 182490 92294
rect 182726 92058 182768 92294
rect 182448 91876 182768 92058
rect 213168 92294 213488 92476
rect 213168 92058 213210 92294
rect 213446 92058 213488 92294
rect 213168 91876 213488 92058
rect 74928 74294 75248 74476
rect 74928 74058 74970 74294
rect 75206 74058 75248 74294
rect 74928 73876 75248 74058
rect 105648 74294 105968 74476
rect 105648 74058 105690 74294
rect 105926 74058 105968 74294
rect 105648 73876 105968 74058
rect 136368 74294 136688 74476
rect 136368 74058 136410 74294
rect 136646 74058 136688 74294
rect 136368 73876 136688 74058
rect 167088 74294 167408 74476
rect 167088 74058 167130 74294
rect 167366 74058 167408 74294
rect 167088 73876 167408 74058
rect 197808 74294 198128 74476
rect 197808 74058 197850 74294
rect 198086 74058 198128 74294
rect 197808 73876 198128 74058
rect 228528 74294 228848 74476
rect 228528 74058 228570 74294
rect 228806 74058 228848 74294
rect 228528 73876 228848 74058
rect 59568 56294 59888 56476
rect 59568 56058 59610 56294
rect 59846 56058 59888 56294
rect 59568 55876 59888 56058
rect 90288 56294 90608 56476
rect 90288 56058 90330 56294
rect 90566 56058 90608 56294
rect 90288 55876 90608 56058
rect 121008 56294 121328 56476
rect 121008 56058 121050 56294
rect 121286 56058 121328 56294
rect 121008 55876 121328 56058
rect 151728 56294 152048 56476
rect 151728 56058 151770 56294
rect 152006 56058 152048 56294
rect 151728 55876 152048 56058
rect 182448 56294 182768 56476
rect 182448 56058 182490 56294
rect 182726 56058 182768 56294
rect 182448 55876 182768 56058
rect 213168 56294 213488 56476
rect 213168 56058 213210 56294
rect 213446 56058 213488 56294
rect 213168 55876 213488 56058
rect 41459 38588 41525 38589
rect 41459 38524 41460 38588
rect 41524 38524 41525 38588
rect 41459 38523 41525 38524
rect 47715 38588 47781 38589
rect 47715 38524 47716 38588
rect 47780 38524 47781 38588
rect 47715 38523 47781 38524
rect 36804 38058 36986 38294
rect 37222 38058 37404 38294
rect 36804 2294 37404 38058
rect 36804 2058 36986 2294
rect 37222 2058 37404 2294
rect 36804 -346 37404 2058
rect 36804 -582 36986 -346
rect 37222 -582 37404 -346
rect 36804 -666 37404 -582
rect 36804 -902 36986 -666
rect 37222 -902 37404 -666
rect 36804 -1894 37404 -902
rect 40504 5994 41104 38000
rect 41462 6221 41522 38523
rect 237422 38453 237482 337315
rect 238504 311994 239104 347758
rect 238504 311758 238686 311994
rect 238922 311758 239104 311994
rect 238504 275994 239104 311758
rect 238504 275758 238686 275994
rect 238922 275758 239104 275994
rect 238504 243568 239104 275758
rect 242204 675694 242804 709082
rect 242204 675458 242386 675694
rect 242622 675458 242804 675694
rect 242204 639694 242804 675458
rect 242204 639458 242386 639694
rect 242622 639458 242804 639694
rect 242204 603694 242804 639458
rect 242204 603458 242386 603694
rect 242622 603458 242804 603694
rect 242204 567694 242804 603458
rect 242204 567458 242386 567694
rect 242622 567458 242804 567694
rect 242204 531694 242804 567458
rect 242204 531458 242386 531694
rect 242622 531458 242804 531694
rect 242204 495694 242804 531458
rect 242204 495458 242386 495694
rect 242622 495458 242804 495694
rect 242204 459694 242804 495458
rect 242204 459458 242386 459694
rect 242622 459458 242804 459694
rect 242204 423694 242804 459458
rect 242204 423458 242386 423694
rect 242622 423458 242804 423694
rect 242204 387694 242804 423458
rect 242204 387458 242386 387694
rect 242622 387458 242804 387694
rect 242204 351694 242804 387458
rect 242204 351458 242386 351694
rect 242622 351458 242804 351694
rect 242204 315694 242804 351458
rect 242204 315458 242386 315694
rect 242622 315458 242804 315694
rect 242204 279694 242804 315458
rect 242204 279458 242386 279694
rect 242622 279458 242804 279694
rect 242204 243694 242804 279458
rect 242204 243458 242386 243694
rect 242622 243458 242804 243694
rect 242204 207694 242804 243458
rect 242204 207458 242386 207694
rect 242622 207458 242804 207694
rect 242204 171694 242804 207458
rect 242204 171458 242386 171694
rect 242622 171458 242804 171694
rect 242204 135694 242804 171458
rect 242204 135458 242386 135694
rect 242622 135458 242804 135694
rect 242204 99694 242804 135458
rect 242204 99458 242386 99694
rect 242622 99458 242804 99694
rect 242204 63694 242804 99458
rect 242204 63458 242386 63694
rect 242622 63458 242804 63694
rect 237419 38452 237485 38453
rect 237419 38388 237420 38452
rect 237484 38388 237485 38452
rect 237419 38387 237485 38388
rect 44204 9694 44804 38000
rect 44204 9458 44386 9694
rect 44622 9458 44804 9694
rect 41459 6220 41525 6221
rect 41459 6156 41460 6220
rect 41524 6156 41525 6220
rect 41459 6155 41525 6156
rect 40504 5758 40686 5994
rect 40922 5758 41104 5994
rect 40504 -2266 41104 5758
rect 40504 -2502 40686 -2266
rect 40922 -2502 41104 -2266
rect 40504 -2586 41104 -2502
rect 40504 -2822 40686 -2586
rect 40922 -2822 41104 -2586
rect 40504 -3814 41104 -2822
rect 44204 -4186 44804 9458
rect 44204 -4422 44386 -4186
rect 44622 -4422 44804 -4186
rect 44204 -4506 44804 -4422
rect 44204 -4742 44386 -4506
rect 44622 -4742 44804 -4506
rect 44204 -5734 44804 -4742
rect 47904 13394 48504 38000
rect 47904 13158 48086 13394
rect 48322 13158 48504 13394
rect 29904 -7302 30086 -7066
rect 30322 -7302 30504 -7066
rect 29904 -7386 30504 -7302
rect 29904 -7622 30086 -7386
rect 30322 -7622 30504 -7386
rect 29904 -7654 30504 -7622
rect 47904 -6106 48504 13158
rect 54804 20294 55404 38000
rect 54804 20058 54986 20294
rect 55222 20058 55404 20294
rect 54804 -1306 55404 20058
rect 54804 -1542 54986 -1306
rect 55222 -1542 55404 -1306
rect 54804 -1626 55404 -1542
rect 54804 -1862 54986 -1626
rect 55222 -1862 55404 -1626
rect 54804 -1894 55404 -1862
rect 58504 23994 59104 38000
rect 58504 23758 58686 23994
rect 58922 23758 59104 23994
rect 58504 -3226 59104 23758
rect 58504 -3462 58686 -3226
rect 58922 -3462 59104 -3226
rect 58504 -3546 59104 -3462
rect 58504 -3782 58686 -3546
rect 58922 -3782 59104 -3546
rect 58504 -3814 59104 -3782
rect 62204 27694 62804 38000
rect 62204 27458 62386 27694
rect 62622 27458 62804 27694
rect 62204 -5146 62804 27458
rect 62204 -5382 62386 -5146
rect 62622 -5382 62804 -5146
rect 62204 -5466 62804 -5382
rect 62204 -5702 62386 -5466
rect 62622 -5702 62804 -5466
rect 62204 -5734 62804 -5702
rect 65904 31394 66504 38000
rect 65904 31158 66086 31394
rect 66322 31158 66504 31394
rect 47904 -6342 48086 -6106
rect 48322 -6342 48504 -6106
rect 47904 -6426 48504 -6342
rect 47904 -6662 48086 -6426
rect 48322 -6662 48504 -6426
rect 47904 -7654 48504 -6662
rect 65904 -7066 66504 31158
rect 72804 2294 73404 38000
rect 72804 2058 72986 2294
rect 73222 2058 73404 2294
rect 72804 -346 73404 2058
rect 72804 -582 72986 -346
rect 73222 -582 73404 -346
rect 72804 -666 73404 -582
rect 72804 -902 72986 -666
rect 73222 -902 73404 -666
rect 72804 -1894 73404 -902
rect 76504 5994 77104 38000
rect 76504 5758 76686 5994
rect 76922 5758 77104 5994
rect 76504 -2266 77104 5758
rect 76504 -2502 76686 -2266
rect 76922 -2502 77104 -2266
rect 76504 -2586 77104 -2502
rect 76504 -2822 76686 -2586
rect 76922 -2822 77104 -2586
rect 76504 -3814 77104 -2822
rect 80204 9694 80804 38000
rect 80204 9458 80386 9694
rect 80622 9458 80804 9694
rect 80204 -4186 80804 9458
rect 80204 -4422 80386 -4186
rect 80622 -4422 80804 -4186
rect 80204 -4506 80804 -4422
rect 80204 -4742 80386 -4506
rect 80622 -4742 80804 -4506
rect 80204 -5734 80804 -4742
rect 83904 13394 84504 38000
rect 83904 13158 84086 13394
rect 84322 13158 84504 13394
rect 65904 -7302 66086 -7066
rect 66322 -7302 66504 -7066
rect 65904 -7386 66504 -7302
rect 65904 -7622 66086 -7386
rect 66322 -7622 66504 -7386
rect 65904 -7654 66504 -7622
rect 83904 -6106 84504 13158
rect 90804 20294 91404 38000
rect 90804 20058 90986 20294
rect 91222 20058 91404 20294
rect 90804 -1306 91404 20058
rect 90804 -1542 90986 -1306
rect 91222 -1542 91404 -1306
rect 90804 -1626 91404 -1542
rect 90804 -1862 90986 -1626
rect 91222 -1862 91404 -1626
rect 90804 -1894 91404 -1862
rect 94504 23994 95104 38000
rect 94504 23758 94686 23994
rect 94922 23758 95104 23994
rect 94504 -3226 95104 23758
rect 94504 -3462 94686 -3226
rect 94922 -3462 95104 -3226
rect 94504 -3546 95104 -3462
rect 94504 -3782 94686 -3546
rect 94922 -3782 95104 -3546
rect 94504 -3814 95104 -3782
rect 98204 27694 98804 38000
rect 98204 27458 98386 27694
rect 98622 27458 98804 27694
rect 98204 -5146 98804 27458
rect 98204 -5382 98386 -5146
rect 98622 -5382 98804 -5146
rect 98204 -5466 98804 -5382
rect 98204 -5702 98386 -5466
rect 98622 -5702 98804 -5466
rect 98204 -5734 98804 -5702
rect 101904 31394 102504 38000
rect 101904 31158 102086 31394
rect 102322 31158 102504 31394
rect 83904 -6342 84086 -6106
rect 84322 -6342 84504 -6106
rect 83904 -6426 84504 -6342
rect 83904 -6662 84086 -6426
rect 84322 -6662 84504 -6426
rect 83904 -7654 84504 -6662
rect 101904 -7066 102504 31158
rect 108804 2294 109404 38000
rect 108804 2058 108986 2294
rect 109222 2058 109404 2294
rect 108804 -346 109404 2058
rect 108804 -582 108986 -346
rect 109222 -582 109404 -346
rect 108804 -666 109404 -582
rect 108804 -902 108986 -666
rect 109222 -902 109404 -666
rect 108804 -1894 109404 -902
rect 112504 5994 113104 38000
rect 112504 5758 112686 5994
rect 112922 5758 113104 5994
rect 112504 -2266 113104 5758
rect 112504 -2502 112686 -2266
rect 112922 -2502 113104 -2266
rect 112504 -2586 113104 -2502
rect 112504 -2822 112686 -2586
rect 112922 -2822 113104 -2586
rect 112504 -3814 113104 -2822
rect 116204 9694 116804 38000
rect 116204 9458 116386 9694
rect 116622 9458 116804 9694
rect 116204 -4186 116804 9458
rect 116204 -4422 116386 -4186
rect 116622 -4422 116804 -4186
rect 116204 -4506 116804 -4422
rect 116204 -4742 116386 -4506
rect 116622 -4742 116804 -4506
rect 116204 -5734 116804 -4742
rect 119904 13394 120504 38000
rect 119904 13158 120086 13394
rect 120322 13158 120504 13394
rect 101904 -7302 102086 -7066
rect 102322 -7302 102504 -7066
rect 101904 -7386 102504 -7302
rect 101904 -7622 102086 -7386
rect 102322 -7622 102504 -7386
rect 101904 -7654 102504 -7622
rect 119904 -6106 120504 13158
rect 126804 20294 127404 38000
rect 126804 20058 126986 20294
rect 127222 20058 127404 20294
rect 126804 -1306 127404 20058
rect 126804 -1542 126986 -1306
rect 127222 -1542 127404 -1306
rect 126804 -1626 127404 -1542
rect 126804 -1862 126986 -1626
rect 127222 -1862 127404 -1626
rect 126804 -1894 127404 -1862
rect 130504 23994 131104 38000
rect 130504 23758 130686 23994
rect 130922 23758 131104 23994
rect 130504 -3226 131104 23758
rect 130504 -3462 130686 -3226
rect 130922 -3462 131104 -3226
rect 130504 -3546 131104 -3462
rect 130504 -3782 130686 -3546
rect 130922 -3782 131104 -3546
rect 130504 -3814 131104 -3782
rect 134204 27694 134804 38000
rect 134204 27458 134386 27694
rect 134622 27458 134804 27694
rect 134204 -5146 134804 27458
rect 134204 -5382 134386 -5146
rect 134622 -5382 134804 -5146
rect 134204 -5466 134804 -5382
rect 134204 -5702 134386 -5466
rect 134622 -5702 134804 -5466
rect 134204 -5734 134804 -5702
rect 137904 31394 138504 38000
rect 137904 31158 138086 31394
rect 138322 31158 138504 31394
rect 119904 -6342 120086 -6106
rect 120322 -6342 120504 -6106
rect 119904 -6426 120504 -6342
rect 119904 -6662 120086 -6426
rect 120322 -6662 120504 -6426
rect 119904 -7654 120504 -6662
rect 137904 -7066 138504 31158
rect 144804 2294 145404 38000
rect 144804 2058 144986 2294
rect 145222 2058 145404 2294
rect 144804 -346 145404 2058
rect 144804 -582 144986 -346
rect 145222 -582 145404 -346
rect 144804 -666 145404 -582
rect 144804 -902 144986 -666
rect 145222 -902 145404 -666
rect 144804 -1894 145404 -902
rect 148504 5994 149104 38000
rect 148504 5758 148686 5994
rect 148922 5758 149104 5994
rect 148504 -2266 149104 5758
rect 148504 -2502 148686 -2266
rect 148922 -2502 149104 -2266
rect 148504 -2586 149104 -2502
rect 148504 -2822 148686 -2586
rect 148922 -2822 149104 -2586
rect 148504 -3814 149104 -2822
rect 152204 9694 152804 38000
rect 152204 9458 152386 9694
rect 152622 9458 152804 9694
rect 152204 -4186 152804 9458
rect 152204 -4422 152386 -4186
rect 152622 -4422 152804 -4186
rect 152204 -4506 152804 -4422
rect 152204 -4742 152386 -4506
rect 152622 -4742 152804 -4506
rect 152204 -5734 152804 -4742
rect 155904 13394 156504 38000
rect 155904 13158 156086 13394
rect 156322 13158 156504 13394
rect 137904 -7302 138086 -7066
rect 138322 -7302 138504 -7066
rect 137904 -7386 138504 -7302
rect 137904 -7622 138086 -7386
rect 138322 -7622 138504 -7386
rect 137904 -7654 138504 -7622
rect 155904 -6106 156504 13158
rect 162804 20294 163404 38000
rect 162804 20058 162986 20294
rect 163222 20058 163404 20294
rect 162804 -1306 163404 20058
rect 162804 -1542 162986 -1306
rect 163222 -1542 163404 -1306
rect 162804 -1626 163404 -1542
rect 162804 -1862 162986 -1626
rect 163222 -1862 163404 -1626
rect 162804 -1894 163404 -1862
rect 166504 23994 167104 38000
rect 166504 23758 166686 23994
rect 166922 23758 167104 23994
rect 166504 -3226 167104 23758
rect 166504 -3462 166686 -3226
rect 166922 -3462 167104 -3226
rect 166504 -3546 167104 -3462
rect 166504 -3782 166686 -3546
rect 166922 -3782 167104 -3546
rect 166504 -3814 167104 -3782
rect 170204 27694 170804 38000
rect 170204 27458 170386 27694
rect 170622 27458 170804 27694
rect 170204 -5146 170804 27458
rect 170204 -5382 170386 -5146
rect 170622 -5382 170804 -5146
rect 170204 -5466 170804 -5382
rect 170204 -5702 170386 -5466
rect 170622 -5702 170804 -5466
rect 170204 -5734 170804 -5702
rect 173904 31394 174504 38000
rect 173904 31158 174086 31394
rect 174322 31158 174504 31394
rect 155904 -6342 156086 -6106
rect 156322 -6342 156504 -6106
rect 155904 -6426 156504 -6342
rect 155904 -6662 156086 -6426
rect 156322 -6662 156504 -6426
rect 155904 -7654 156504 -6662
rect 173904 -7066 174504 31158
rect 180804 2294 181404 38000
rect 180804 2058 180986 2294
rect 181222 2058 181404 2294
rect 180804 -346 181404 2058
rect 180804 -582 180986 -346
rect 181222 -582 181404 -346
rect 180804 -666 181404 -582
rect 180804 -902 180986 -666
rect 181222 -902 181404 -666
rect 180804 -1894 181404 -902
rect 184504 5994 185104 38000
rect 184504 5758 184686 5994
rect 184922 5758 185104 5994
rect 184504 -2266 185104 5758
rect 184504 -2502 184686 -2266
rect 184922 -2502 185104 -2266
rect 184504 -2586 185104 -2502
rect 184504 -2822 184686 -2586
rect 184922 -2822 185104 -2586
rect 184504 -3814 185104 -2822
rect 188204 9694 188804 38000
rect 188204 9458 188386 9694
rect 188622 9458 188804 9694
rect 188204 -4186 188804 9458
rect 188204 -4422 188386 -4186
rect 188622 -4422 188804 -4186
rect 188204 -4506 188804 -4422
rect 188204 -4742 188386 -4506
rect 188622 -4742 188804 -4506
rect 188204 -5734 188804 -4742
rect 191904 13394 192504 38000
rect 191904 13158 192086 13394
rect 192322 13158 192504 13394
rect 173904 -7302 174086 -7066
rect 174322 -7302 174504 -7066
rect 173904 -7386 174504 -7302
rect 173904 -7622 174086 -7386
rect 174322 -7622 174504 -7386
rect 173904 -7654 174504 -7622
rect 191904 -6106 192504 13158
rect 198804 20294 199404 38000
rect 198804 20058 198986 20294
rect 199222 20058 199404 20294
rect 198804 -1306 199404 20058
rect 198804 -1542 198986 -1306
rect 199222 -1542 199404 -1306
rect 198804 -1626 199404 -1542
rect 198804 -1862 198986 -1626
rect 199222 -1862 199404 -1626
rect 198804 -1894 199404 -1862
rect 202504 23994 203104 38000
rect 202504 23758 202686 23994
rect 202922 23758 203104 23994
rect 202504 -3226 203104 23758
rect 202504 -3462 202686 -3226
rect 202922 -3462 203104 -3226
rect 202504 -3546 203104 -3462
rect 202504 -3782 202686 -3546
rect 202922 -3782 203104 -3546
rect 202504 -3814 203104 -3782
rect 206204 27694 206804 38000
rect 206204 27458 206386 27694
rect 206622 27458 206804 27694
rect 206204 -5146 206804 27458
rect 206204 -5382 206386 -5146
rect 206622 -5382 206804 -5146
rect 206204 -5466 206804 -5382
rect 206204 -5702 206386 -5466
rect 206622 -5702 206804 -5466
rect 206204 -5734 206804 -5702
rect 209904 31394 210504 38000
rect 209904 31158 210086 31394
rect 210322 31158 210504 31394
rect 191904 -6342 192086 -6106
rect 192322 -6342 192504 -6106
rect 191904 -6426 192504 -6342
rect 191904 -6662 192086 -6426
rect 192322 -6662 192504 -6426
rect 191904 -7654 192504 -6662
rect 209904 -7066 210504 31158
rect 216804 2294 217404 38000
rect 216804 2058 216986 2294
rect 217222 2058 217404 2294
rect 216804 -346 217404 2058
rect 216804 -582 216986 -346
rect 217222 -582 217404 -346
rect 216804 -666 217404 -582
rect 216804 -902 216986 -666
rect 217222 -902 217404 -666
rect 216804 -1894 217404 -902
rect 220504 5994 221104 38000
rect 220504 5758 220686 5994
rect 220922 5758 221104 5994
rect 220504 -2266 221104 5758
rect 220504 -2502 220686 -2266
rect 220922 -2502 221104 -2266
rect 220504 -2586 221104 -2502
rect 220504 -2822 220686 -2586
rect 220922 -2822 221104 -2586
rect 220504 -3814 221104 -2822
rect 224204 9694 224804 38000
rect 224204 9458 224386 9694
rect 224622 9458 224804 9694
rect 224204 -4186 224804 9458
rect 224204 -4422 224386 -4186
rect 224622 -4422 224804 -4186
rect 224204 -4506 224804 -4422
rect 224204 -4742 224386 -4506
rect 224622 -4742 224804 -4506
rect 224204 -5734 224804 -4742
rect 227904 13394 228504 38000
rect 227904 13158 228086 13394
rect 228322 13158 228504 13394
rect 209904 -7302 210086 -7066
rect 210322 -7302 210504 -7066
rect 209904 -7386 210504 -7302
rect 209904 -7622 210086 -7386
rect 210322 -7622 210504 -7386
rect 209904 -7654 210504 -7622
rect 227904 -6106 228504 13158
rect 234804 20294 235404 38000
rect 234804 20058 234986 20294
rect 235222 20058 235404 20294
rect 234804 -1306 235404 20058
rect 234804 -1542 234986 -1306
rect 235222 -1542 235404 -1306
rect 234804 -1626 235404 -1542
rect 234804 -1862 234986 -1626
rect 235222 -1862 235404 -1626
rect 234804 -1894 235404 -1862
rect 238504 23994 239104 38000
rect 238504 23758 238686 23994
rect 238922 23758 239104 23994
rect 238504 -3226 239104 23758
rect 238504 -3462 238686 -3226
rect 238922 -3462 239104 -3226
rect 238504 -3546 239104 -3462
rect 238504 -3782 238686 -3546
rect 238922 -3782 239104 -3546
rect 238504 -3814 239104 -3782
rect 242204 27694 242804 63458
rect 242204 27458 242386 27694
rect 242622 27458 242804 27694
rect 242204 -5146 242804 27458
rect 242204 -5382 242386 -5146
rect 242622 -5382 242804 -5146
rect 242204 -5466 242804 -5382
rect 242204 -5702 242386 -5466
rect 242622 -5702 242804 -5466
rect 242204 -5734 242804 -5702
rect 245904 679394 246504 711002
rect 263904 710598 264504 711590
rect 263904 710362 264086 710598
rect 264322 710362 264504 710598
rect 263904 710278 264504 710362
rect 263904 710042 264086 710278
rect 264322 710042 264504 710278
rect 260204 708678 260804 709670
rect 260204 708442 260386 708678
rect 260622 708442 260804 708678
rect 260204 708358 260804 708442
rect 260204 708122 260386 708358
rect 260622 708122 260804 708358
rect 256504 706758 257104 707750
rect 256504 706522 256686 706758
rect 256922 706522 257104 706758
rect 256504 706438 257104 706522
rect 256504 706202 256686 706438
rect 256922 706202 257104 706438
rect 245904 679158 246086 679394
rect 246322 679158 246504 679394
rect 245904 643394 246504 679158
rect 245904 643158 246086 643394
rect 246322 643158 246504 643394
rect 245904 607394 246504 643158
rect 245904 607158 246086 607394
rect 246322 607158 246504 607394
rect 245904 571394 246504 607158
rect 245904 571158 246086 571394
rect 246322 571158 246504 571394
rect 245904 535394 246504 571158
rect 245904 535158 246086 535394
rect 246322 535158 246504 535394
rect 245904 499394 246504 535158
rect 245904 499158 246086 499394
rect 246322 499158 246504 499394
rect 245904 463394 246504 499158
rect 245904 463158 246086 463394
rect 246322 463158 246504 463394
rect 245904 427394 246504 463158
rect 245904 427158 246086 427394
rect 246322 427158 246504 427394
rect 245904 391394 246504 427158
rect 245904 391158 246086 391394
rect 246322 391158 246504 391394
rect 245904 355394 246504 391158
rect 245904 355158 246086 355394
rect 246322 355158 246504 355394
rect 245904 319394 246504 355158
rect 245904 319158 246086 319394
rect 246322 319158 246504 319394
rect 245904 283394 246504 319158
rect 245904 283158 246086 283394
rect 246322 283158 246504 283394
rect 245904 247394 246504 283158
rect 245904 247158 246086 247394
rect 246322 247158 246504 247394
rect 245904 211394 246504 247158
rect 245904 211158 246086 211394
rect 246322 211158 246504 211394
rect 245904 175394 246504 211158
rect 245904 175158 246086 175394
rect 246322 175158 246504 175394
rect 245904 139394 246504 175158
rect 245904 139158 246086 139394
rect 246322 139158 246504 139394
rect 245904 103394 246504 139158
rect 245904 103158 246086 103394
rect 246322 103158 246504 103394
rect 245904 67394 246504 103158
rect 245904 67158 246086 67394
rect 246322 67158 246504 67394
rect 245904 31394 246504 67158
rect 245904 31158 246086 31394
rect 246322 31158 246504 31394
rect 227904 -6342 228086 -6106
rect 228322 -6342 228504 -6106
rect 227904 -6426 228504 -6342
rect 227904 -6662 228086 -6426
rect 228322 -6662 228504 -6426
rect 227904 -7654 228504 -6662
rect 245904 -7066 246504 31158
rect 252804 704838 253404 705830
rect 252804 704602 252986 704838
rect 253222 704602 253404 704838
rect 252804 704518 253404 704602
rect 252804 704282 252986 704518
rect 253222 704282 253404 704518
rect 252804 686294 253404 704282
rect 252804 686058 252986 686294
rect 253222 686058 253404 686294
rect 252804 650294 253404 686058
rect 252804 650058 252986 650294
rect 253222 650058 253404 650294
rect 252804 614294 253404 650058
rect 252804 614058 252986 614294
rect 253222 614058 253404 614294
rect 252804 578294 253404 614058
rect 252804 578058 252986 578294
rect 253222 578058 253404 578294
rect 252804 542294 253404 578058
rect 252804 542058 252986 542294
rect 253222 542058 253404 542294
rect 252804 506294 253404 542058
rect 252804 506058 252986 506294
rect 253222 506058 253404 506294
rect 252804 470294 253404 506058
rect 252804 470058 252986 470294
rect 253222 470058 253404 470294
rect 252804 434294 253404 470058
rect 252804 434058 252986 434294
rect 253222 434058 253404 434294
rect 252804 398294 253404 434058
rect 252804 398058 252986 398294
rect 253222 398058 253404 398294
rect 252804 362294 253404 398058
rect 252804 362058 252986 362294
rect 253222 362058 253404 362294
rect 252804 326294 253404 362058
rect 252804 326058 252986 326294
rect 253222 326058 253404 326294
rect 252804 290294 253404 326058
rect 252804 290058 252986 290294
rect 253222 290058 253404 290294
rect 252804 254294 253404 290058
rect 252804 254058 252986 254294
rect 253222 254058 253404 254294
rect 252804 218294 253404 254058
rect 252804 218058 252986 218294
rect 253222 218058 253404 218294
rect 252804 182294 253404 218058
rect 252804 182058 252986 182294
rect 253222 182058 253404 182294
rect 252804 146294 253404 182058
rect 252804 146058 252986 146294
rect 253222 146058 253404 146294
rect 252804 110294 253404 146058
rect 252804 110058 252986 110294
rect 253222 110058 253404 110294
rect 252804 74294 253404 110058
rect 252804 74058 252986 74294
rect 253222 74058 253404 74294
rect 252804 38294 253404 74058
rect 252804 38058 252986 38294
rect 253222 38058 253404 38294
rect 252804 2294 253404 38058
rect 252804 2058 252986 2294
rect 253222 2058 253404 2294
rect 252804 -346 253404 2058
rect 252804 -582 252986 -346
rect 253222 -582 253404 -346
rect 252804 -666 253404 -582
rect 252804 -902 252986 -666
rect 253222 -902 253404 -666
rect 252804 -1894 253404 -902
rect 256504 689994 257104 706202
rect 256504 689758 256686 689994
rect 256922 689758 257104 689994
rect 256504 653994 257104 689758
rect 256504 653758 256686 653994
rect 256922 653758 257104 653994
rect 256504 617994 257104 653758
rect 256504 617758 256686 617994
rect 256922 617758 257104 617994
rect 256504 581994 257104 617758
rect 256504 581758 256686 581994
rect 256922 581758 257104 581994
rect 256504 545994 257104 581758
rect 256504 545758 256686 545994
rect 256922 545758 257104 545994
rect 256504 509994 257104 545758
rect 256504 509758 256686 509994
rect 256922 509758 257104 509994
rect 256504 473994 257104 509758
rect 256504 473758 256686 473994
rect 256922 473758 257104 473994
rect 256504 437994 257104 473758
rect 256504 437758 256686 437994
rect 256922 437758 257104 437994
rect 256504 401994 257104 437758
rect 256504 401758 256686 401994
rect 256922 401758 257104 401994
rect 256504 365994 257104 401758
rect 256504 365758 256686 365994
rect 256922 365758 257104 365994
rect 256504 329994 257104 365758
rect 256504 329758 256686 329994
rect 256922 329758 257104 329994
rect 256504 293994 257104 329758
rect 256504 293758 256686 293994
rect 256922 293758 257104 293994
rect 256504 257994 257104 293758
rect 256504 257758 256686 257994
rect 256922 257758 257104 257994
rect 256504 221994 257104 257758
rect 256504 221758 256686 221994
rect 256922 221758 257104 221994
rect 256504 185994 257104 221758
rect 256504 185758 256686 185994
rect 256922 185758 257104 185994
rect 256504 149994 257104 185758
rect 256504 149758 256686 149994
rect 256922 149758 257104 149994
rect 256504 113994 257104 149758
rect 256504 113758 256686 113994
rect 256922 113758 257104 113994
rect 256504 77994 257104 113758
rect 256504 77758 256686 77994
rect 256922 77758 257104 77994
rect 256504 41994 257104 77758
rect 256504 41758 256686 41994
rect 256922 41758 257104 41994
rect 256504 5994 257104 41758
rect 256504 5758 256686 5994
rect 256922 5758 257104 5994
rect 256504 -2266 257104 5758
rect 256504 -2502 256686 -2266
rect 256922 -2502 257104 -2266
rect 256504 -2586 257104 -2502
rect 256504 -2822 256686 -2586
rect 256922 -2822 257104 -2586
rect 256504 -3814 257104 -2822
rect 260204 693694 260804 708122
rect 260204 693458 260386 693694
rect 260622 693458 260804 693694
rect 260204 657694 260804 693458
rect 260204 657458 260386 657694
rect 260622 657458 260804 657694
rect 260204 621694 260804 657458
rect 260204 621458 260386 621694
rect 260622 621458 260804 621694
rect 260204 585694 260804 621458
rect 260204 585458 260386 585694
rect 260622 585458 260804 585694
rect 260204 549694 260804 585458
rect 260204 549458 260386 549694
rect 260622 549458 260804 549694
rect 260204 513694 260804 549458
rect 260204 513458 260386 513694
rect 260622 513458 260804 513694
rect 260204 477694 260804 513458
rect 260204 477458 260386 477694
rect 260622 477458 260804 477694
rect 260204 441694 260804 477458
rect 260204 441458 260386 441694
rect 260622 441458 260804 441694
rect 260204 405694 260804 441458
rect 260204 405458 260386 405694
rect 260622 405458 260804 405694
rect 260204 369694 260804 405458
rect 260204 369458 260386 369694
rect 260622 369458 260804 369694
rect 260204 333694 260804 369458
rect 260204 333458 260386 333694
rect 260622 333458 260804 333694
rect 260204 297694 260804 333458
rect 260204 297458 260386 297694
rect 260622 297458 260804 297694
rect 260204 261694 260804 297458
rect 260204 261458 260386 261694
rect 260622 261458 260804 261694
rect 260204 225694 260804 261458
rect 260204 225458 260386 225694
rect 260622 225458 260804 225694
rect 260204 189694 260804 225458
rect 260204 189458 260386 189694
rect 260622 189458 260804 189694
rect 260204 153694 260804 189458
rect 260204 153458 260386 153694
rect 260622 153458 260804 153694
rect 260204 117694 260804 153458
rect 260204 117458 260386 117694
rect 260622 117458 260804 117694
rect 260204 81694 260804 117458
rect 260204 81458 260386 81694
rect 260622 81458 260804 81694
rect 260204 45694 260804 81458
rect 260204 45458 260386 45694
rect 260622 45458 260804 45694
rect 260204 9694 260804 45458
rect 260204 9458 260386 9694
rect 260622 9458 260804 9694
rect 260204 -4186 260804 9458
rect 260204 -4422 260386 -4186
rect 260622 -4422 260804 -4186
rect 260204 -4506 260804 -4422
rect 260204 -4742 260386 -4506
rect 260622 -4742 260804 -4506
rect 260204 -5734 260804 -4742
rect 263904 697394 264504 710042
rect 281904 711558 282504 711590
rect 281904 711322 282086 711558
rect 282322 711322 282504 711558
rect 281904 711238 282504 711322
rect 281904 711002 282086 711238
rect 282322 711002 282504 711238
rect 278204 709638 278804 709670
rect 278204 709402 278386 709638
rect 278622 709402 278804 709638
rect 278204 709318 278804 709402
rect 278204 709082 278386 709318
rect 278622 709082 278804 709318
rect 274504 707718 275104 707750
rect 274504 707482 274686 707718
rect 274922 707482 275104 707718
rect 274504 707398 275104 707482
rect 274504 707162 274686 707398
rect 274922 707162 275104 707398
rect 263904 697158 264086 697394
rect 264322 697158 264504 697394
rect 263904 661394 264504 697158
rect 263904 661158 264086 661394
rect 264322 661158 264504 661394
rect 263904 625394 264504 661158
rect 263904 625158 264086 625394
rect 264322 625158 264504 625394
rect 263904 589394 264504 625158
rect 263904 589158 264086 589394
rect 264322 589158 264504 589394
rect 263904 553394 264504 589158
rect 263904 553158 264086 553394
rect 264322 553158 264504 553394
rect 263904 517394 264504 553158
rect 263904 517158 264086 517394
rect 264322 517158 264504 517394
rect 263904 481394 264504 517158
rect 263904 481158 264086 481394
rect 264322 481158 264504 481394
rect 263904 445394 264504 481158
rect 263904 445158 264086 445394
rect 264322 445158 264504 445394
rect 263904 409394 264504 445158
rect 263904 409158 264086 409394
rect 264322 409158 264504 409394
rect 263904 373394 264504 409158
rect 263904 373158 264086 373394
rect 264322 373158 264504 373394
rect 263904 337394 264504 373158
rect 263904 337158 264086 337394
rect 264322 337158 264504 337394
rect 263904 301394 264504 337158
rect 263904 301158 264086 301394
rect 264322 301158 264504 301394
rect 263904 265394 264504 301158
rect 263904 265158 264086 265394
rect 264322 265158 264504 265394
rect 263904 229394 264504 265158
rect 263904 229158 264086 229394
rect 264322 229158 264504 229394
rect 263904 193394 264504 229158
rect 263904 193158 264086 193394
rect 264322 193158 264504 193394
rect 263904 157394 264504 193158
rect 263904 157158 264086 157394
rect 264322 157158 264504 157394
rect 263904 121394 264504 157158
rect 263904 121158 264086 121394
rect 264322 121158 264504 121394
rect 263904 85394 264504 121158
rect 263904 85158 264086 85394
rect 264322 85158 264504 85394
rect 263904 49394 264504 85158
rect 263904 49158 264086 49394
rect 264322 49158 264504 49394
rect 263904 13394 264504 49158
rect 263904 13158 264086 13394
rect 264322 13158 264504 13394
rect 245904 -7302 246086 -7066
rect 246322 -7302 246504 -7066
rect 245904 -7386 246504 -7302
rect 245904 -7622 246086 -7386
rect 246322 -7622 246504 -7386
rect 245904 -7654 246504 -7622
rect 263904 -6106 264504 13158
rect 270804 705798 271404 705830
rect 270804 705562 270986 705798
rect 271222 705562 271404 705798
rect 270804 705478 271404 705562
rect 270804 705242 270986 705478
rect 271222 705242 271404 705478
rect 270804 668294 271404 705242
rect 270804 668058 270986 668294
rect 271222 668058 271404 668294
rect 270804 632294 271404 668058
rect 270804 632058 270986 632294
rect 271222 632058 271404 632294
rect 270804 596294 271404 632058
rect 270804 596058 270986 596294
rect 271222 596058 271404 596294
rect 270804 560294 271404 596058
rect 270804 560058 270986 560294
rect 271222 560058 271404 560294
rect 270804 524294 271404 560058
rect 270804 524058 270986 524294
rect 271222 524058 271404 524294
rect 270804 488294 271404 524058
rect 270804 488058 270986 488294
rect 271222 488058 271404 488294
rect 270804 452294 271404 488058
rect 270804 452058 270986 452294
rect 271222 452058 271404 452294
rect 270804 416294 271404 452058
rect 270804 416058 270986 416294
rect 271222 416058 271404 416294
rect 270804 380294 271404 416058
rect 270804 380058 270986 380294
rect 271222 380058 271404 380294
rect 270804 344294 271404 380058
rect 270804 344058 270986 344294
rect 271222 344058 271404 344294
rect 270804 308294 271404 344058
rect 270804 308058 270986 308294
rect 271222 308058 271404 308294
rect 270804 272294 271404 308058
rect 270804 272058 270986 272294
rect 271222 272058 271404 272294
rect 270804 236294 271404 272058
rect 270804 236058 270986 236294
rect 271222 236058 271404 236294
rect 270804 200294 271404 236058
rect 270804 200058 270986 200294
rect 271222 200058 271404 200294
rect 270804 164294 271404 200058
rect 270804 164058 270986 164294
rect 271222 164058 271404 164294
rect 270804 128294 271404 164058
rect 270804 128058 270986 128294
rect 271222 128058 271404 128294
rect 270804 92294 271404 128058
rect 270804 92058 270986 92294
rect 271222 92058 271404 92294
rect 270804 56294 271404 92058
rect 270804 56058 270986 56294
rect 271222 56058 271404 56294
rect 270804 20294 271404 56058
rect 270804 20058 270986 20294
rect 271222 20058 271404 20294
rect 270804 -1306 271404 20058
rect 270804 -1542 270986 -1306
rect 271222 -1542 271404 -1306
rect 270804 -1626 271404 -1542
rect 270804 -1862 270986 -1626
rect 271222 -1862 271404 -1626
rect 270804 -1894 271404 -1862
rect 274504 671994 275104 707162
rect 274504 671758 274686 671994
rect 274922 671758 275104 671994
rect 274504 635994 275104 671758
rect 274504 635758 274686 635994
rect 274922 635758 275104 635994
rect 274504 599994 275104 635758
rect 274504 599758 274686 599994
rect 274922 599758 275104 599994
rect 274504 563994 275104 599758
rect 274504 563758 274686 563994
rect 274922 563758 275104 563994
rect 274504 527994 275104 563758
rect 274504 527758 274686 527994
rect 274922 527758 275104 527994
rect 274504 491994 275104 527758
rect 274504 491758 274686 491994
rect 274922 491758 275104 491994
rect 274504 455994 275104 491758
rect 274504 455758 274686 455994
rect 274922 455758 275104 455994
rect 274504 419994 275104 455758
rect 274504 419758 274686 419994
rect 274922 419758 275104 419994
rect 274504 383994 275104 419758
rect 274504 383758 274686 383994
rect 274922 383758 275104 383994
rect 274504 347994 275104 383758
rect 274504 347758 274686 347994
rect 274922 347758 275104 347994
rect 274504 311994 275104 347758
rect 274504 311758 274686 311994
rect 274922 311758 275104 311994
rect 274504 275994 275104 311758
rect 274504 275758 274686 275994
rect 274922 275758 275104 275994
rect 274504 239994 275104 275758
rect 274504 239758 274686 239994
rect 274922 239758 275104 239994
rect 274504 203994 275104 239758
rect 274504 203758 274686 203994
rect 274922 203758 275104 203994
rect 274504 167994 275104 203758
rect 274504 167758 274686 167994
rect 274922 167758 275104 167994
rect 274504 131994 275104 167758
rect 274504 131758 274686 131994
rect 274922 131758 275104 131994
rect 274504 95994 275104 131758
rect 274504 95758 274686 95994
rect 274922 95758 275104 95994
rect 274504 59994 275104 95758
rect 274504 59758 274686 59994
rect 274922 59758 275104 59994
rect 274504 23994 275104 59758
rect 274504 23758 274686 23994
rect 274922 23758 275104 23994
rect 274504 -3226 275104 23758
rect 274504 -3462 274686 -3226
rect 274922 -3462 275104 -3226
rect 274504 -3546 275104 -3462
rect 274504 -3782 274686 -3546
rect 274922 -3782 275104 -3546
rect 274504 -3814 275104 -3782
rect 278204 675694 278804 709082
rect 278204 675458 278386 675694
rect 278622 675458 278804 675694
rect 278204 639694 278804 675458
rect 278204 639458 278386 639694
rect 278622 639458 278804 639694
rect 278204 603694 278804 639458
rect 278204 603458 278386 603694
rect 278622 603458 278804 603694
rect 278204 567694 278804 603458
rect 278204 567458 278386 567694
rect 278622 567458 278804 567694
rect 278204 531694 278804 567458
rect 278204 531458 278386 531694
rect 278622 531458 278804 531694
rect 278204 495694 278804 531458
rect 278204 495458 278386 495694
rect 278622 495458 278804 495694
rect 278204 459694 278804 495458
rect 278204 459458 278386 459694
rect 278622 459458 278804 459694
rect 278204 423694 278804 459458
rect 278204 423458 278386 423694
rect 278622 423458 278804 423694
rect 278204 387694 278804 423458
rect 278204 387458 278386 387694
rect 278622 387458 278804 387694
rect 278204 351694 278804 387458
rect 278204 351458 278386 351694
rect 278622 351458 278804 351694
rect 278204 315694 278804 351458
rect 278204 315458 278386 315694
rect 278622 315458 278804 315694
rect 278204 279694 278804 315458
rect 278204 279458 278386 279694
rect 278622 279458 278804 279694
rect 278204 243694 278804 279458
rect 278204 243458 278386 243694
rect 278622 243458 278804 243694
rect 278204 207694 278804 243458
rect 278204 207458 278386 207694
rect 278622 207458 278804 207694
rect 278204 171694 278804 207458
rect 278204 171458 278386 171694
rect 278622 171458 278804 171694
rect 278204 135694 278804 171458
rect 278204 135458 278386 135694
rect 278622 135458 278804 135694
rect 278204 99694 278804 135458
rect 278204 99458 278386 99694
rect 278622 99458 278804 99694
rect 278204 63694 278804 99458
rect 278204 63458 278386 63694
rect 278622 63458 278804 63694
rect 278204 27694 278804 63458
rect 278204 27458 278386 27694
rect 278622 27458 278804 27694
rect 278204 -5146 278804 27458
rect 278204 -5382 278386 -5146
rect 278622 -5382 278804 -5146
rect 278204 -5466 278804 -5382
rect 278204 -5702 278386 -5466
rect 278622 -5702 278804 -5466
rect 278204 -5734 278804 -5702
rect 281904 679394 282504 711002
rect 299904 710598 300504 711590
rect 299904 710362 300086 710598
rect 300322 710362 300504 710598
rect 299904 710278 300504 710362
rect 299904 710042 300086 710278
rect 300322 710042 300504 710278
rect 296204 708678 296804 709670
rect 296204 708442 296386 708678
rect 296622 708442 296804 708678
rect 296204 708358 296804 708442
rect 296204 708122 296386 708358
rect 296622 708122 296804 708358
rect 292504 706758 293104 707750
rect 292504 706522 292686 706758
rect 292922 706522 293104 706758
rect 292504 706438 293104 706522
rect 292504 706202 292686 706438
rect 292922 706202 293104 706438
rect 281904 679158 282086 679394
rect 282322 679158 282504 679394
rect 281904 643394 282504 679158
rect 281904 643158 282086 643394
rect 282322 643158 282504 643394
rect 281904 607394 282504 643158
rect 281904 607158 282086 607394
rect 282322 607158 282504 607394
rect 281904 571394 282504 607158
rect 281904 571158 282086 571394
rect 282322 571158 282504 571394
rect 281904 535394 282504 571158
rect 281904 535158 282086 535394
rect 282322 535158 282504 535394
rect 281904 499394 282504 535158
rect 281904 499158 282086 499394
rect 282322 499158 282504 499394
rect 281904 463394 282504 499158
rect 281904 463158 282086 463394
rect 282322 463158 282504 463394
rect 281904 427394 282504 463158
rect 281904 427158 282086 427394
rect 282322 427158 282504 427394
rect 281904 391394 282504 427158
rect 281904 391158 282086 391394
rect 282322 391158 282504 391394
rect 281904 355394 282504 391158
rect 281904 355158 282086 355394
rect 282322 355158 282504 355394
rect 281904 319394 282504 355158
rect 281904 319158 282086 319394
rect 282322 319158 282504 319394
rect 281904 283394 282504 319158
rect 281904 283158 282086 283394
rect 282322 283158 282504 283394
rect 281904 247394 282504 283158
rect 281904 247158 282086 247394
rect 282322 247158 282504 247394
rect 281904 211394 282504 247158
rect 281904 211158 282086 211394
rect 282322 211158 282504 211394
rect 281904 175394 282504 211158
rect 281904 175158 282086 175394
rect 282322 175158 282504 175394
rect 281904 139394 282504 175158
rect 281904 139158 282086 139394
rect 282322 139158 282504 139394
rect 281904 103394 282504 139158
rect 281904 103158 282086 103394
rect 282322 103158 282504 103394
rect 281904 67394 282504 103158
rect 281904 67158 282086 67394
rect 282322 67158 282504 67394
rect 281904 31394 282504 67158
rect 281904 31158 282086 31394
rect 282322 31158 282504 31394
rect 263904 -6342 264086 -6106
rect 264322 -6342 264504 -6106
rect 263904 -6426 264504 -6342
rect 263904 -6662 264086 -6426
rect 264322 -6662 264504 -6426
rect 263904 -7654 264504 -6662
rect 281904 -7066 282504 31158
rect 288804 704838 289404 705830
rect 288804 704602 288986 704838
rect 289222 704602 289404 704838
rect 288804 704518 289404 704602
rect 288804 704282 288986 704518
rect 289222 704282 289404 704518
rect 288804 686294 289404 704282
rect 288804 686058 288986 686294
rect 289222 686058 289404 686294
rect 288804 650294 289404 686058
rect 288804 650058 288986 650294
rect 289222 650058 289404 650294
rect 288804 614294 289404 650058
rect 288804 614058 288986 614294
rect 289222 614058 289404 614294
rect 288804 578294 289404 614058
rect 288804 578058 288986 578294
rect 289222 578058 289404 578294
rect 288804 542294 289404 578058
rect 288804 542058 288986 542294
rect 289222 542058 289404 542294
rect 288804 506294 289404 542058
rect 288804 506058 288986 506294
rect 289222 506058 289404 506294
rect 288804 470294 289404 506058
rect 288804 470058 288986 470294
rect 289222 470058 289404 470294
rect 288804 434294 289404 470058
rect 288804 434058 288986 434294
rect 289222 434058 289404 434294
rect 288804 398294 289404 434058
rect 288804 398058 288986 398294
rect 289222 398058 289404 398294
rect 288804 362294 289404 398058
rect 288804 362058 288986 362294
rect 289222 362058 289404 362294
rect 288804 326294 289404 362058
rect 288804 326058 288986 326294
rect 289222 326058 289404 326294
rect 288804 290294 289404 326058
rect 288804 290058 288986 290294
rect 289222 290058 289404 290294
rect 288804 254294 289404 290058
rect 288804 254058 288986 254294
rect 289222 254058 289404 254294
rect 288804 218294 289404 254058
rect 288804 218058 288986 218294
rect 289222 218058 289404 218294
rect 288804 182294 289404 218058
rect 288804 182058 288986 182294
rect 289222 182058 289404 182294
rect 288804 146294 289404 182058
rect 288804 146058 288986 146294
rect 289222 146058 289404 146294
rect 288804 110294 289404 146058
rect 288804 110058 288986 110294
rect 289222 110058 289404 110294
rect 288804 74294 289404 110058
rect 288804 74058 288986 74294
rect 289222 74058 289404 74294
rect 288804 38294 289404 74058
rect 288804 38058 288986 38294
rect 289222 38058 289404 38294
rect 288804 2294 289404 38058
rect 288804 2058 288986 2294
rect 289222 2058 289404 2294
rect 288804 -346 289404 2058
rect 288804 -582 288986 -346
rect 289222 -582 289404 -346
rect 288804 -666 289404 -582
rect 288804 -902 288986 -666
rect 289222 -902 289404 -666
rect 288804 -1894 289404 -902
rect 292504 689994 293104 706202
rect 292504 689758 292686 689994
rect 292922 689758 293104 689994
rect 292504 653994 293104 689758
rect 292504 653758 292686 653994
rect 292922 653758 293104 653994
rect 292504 617994 293104 653758
rect 292504 617758 292686 617994
rect 292922 617758 293104 617994
rect 292504 581994 293104 617758
rect 292504 581758 292686 581994
rect 292922 581758 293104 581994
rect 292504 545994 293104 581758
rect 292504 545758 292686 545994
rect 292922 545758 293104 545994
rect 292504 509994 293104 545758
rect 292504 509758 292686 509994
rect 292922 509758 293104 509994
rect 292504 473994 293104 509758
rect 292504 473758 292686 473994
rect 292922 473758 293104 473994
rect 292504 437994 293104 473758
rect 292504 437758 292686 437994
rect 292922 437758 293104 437994
rect 292504 401994 293104 437758
rect 292504 401758 292686 401994
rect 292922 401758 293104 401994
rect 292504 365994 293104 401758
rect 292504 365758 292686 365994
rect 292922 365758 293104 365994
rect 292504 329994 293104 365758
rect 292504 329758 292686 329994
rect 292922 329758 293104 329994
rect 292504 293994 293104 329758
rect 292504 293758 292686 293994
rect 292922 293758 293104 293994
rect 292504 257994 293104 293758
rect 292504 257758 292686 257994
rect 292922 257758 293104 257994
rect 292504 221994 293104 257758
rect 292504 221758 292686 221994
rect 292922 221758 293104 221994
rect 292504 185994 293104 221758
rect 292504 185758 292686 185994
rect 292922 185758 293104 185994
rect 292504 149994 293104 185758
rect 292504 149758 292686 149994
rect 292922 149758 293104 149994
rect 292504 113994 293104 149758
rect 292504 113758 292686 113994
rect 292922 113758 293104 113994
rect 292504 77994 293104 113758
rect 292504 77758 292686 77994
rect 292922 77758 293104 77994
rect 292504 41994 293104 77758
rect 292504 41758 292686 41994
rect 292922 41758 293104 41994
rect 292504 5994 293104 41758
rect 292504 5758 292686 5994
rect 292922 5758 293104 5994
rect 292504 -2266 293104 5758
rect 292504 -2502 292686 -2266
rect 292922 -2502 293104 -2266
rect 292504 -2586 293104 -2502
rect 292504 -2822 292686 -2586
rect 292922 -2822 293104 -2586
rect 292504 -3814 293104 -2822
rect 296204 693694 296804 708122
rect 296204 693458 296386 693694
rect 296622 693458 296804 693694
rect 296204 657694 296804 693458
rect 296204 657458 296386 657694
rect 296622 657458 296804 657694
rect 296204 621694 296804 657458
rect 296204 621458 296386 621694
rect 296622 621458 296804 621694
rect 296204 585694 296804 621458
rect 296204 585458 296386 585694
rect 296622 585458 296804 585694
rect 296204 549694 296804 585458
rect 296204 549458 296386 549694
rect 296622 549458 296804 549694
rect 296204 513694 296804 549458
rect 296204 513458 296386 513694
rect 296622 513458 296804 513694
rect 296204 477694 296804 513458
rect 296204 477458 296386 477694
rect 296622 477458 296804 477694
rect 296204 441694 296804 477458
rect 296204 441458 296386 441694
rect 296622 441458 296804 441694
rect 296204 405694 296804 441458
rect 296204 405458 296386 405694
rect 296622 405458 296804 405694
rect 296204 369694 296804 405458
rect 296204 369458 296386 369694
rect 296622 369458 296804 369694
rect 296204 333694 296804 369458
rect 296204 333458 296386 333694
rect 296622 333458 296804 333694
rect 296204 297694 296804 333458
rect 296204 297458 296386 297694
rect 296622 297458 296804 297694
rect 296204 261694 296804 297458
rect 296204 261458 296386 261694
rect 296622 261458 296804 261694
rect 296204 225694 296804 261458
rect 296204 225458 296386 225694
rect 296622 225458 296804 225694
rect 296204 189694 296804 225458
rect 296204 189458 296386 189694
rect 296622 189458 296804 189694
rect 296204 153694 296804 189458
rect 296204 153458 296386 153694
rect 296622 153458 296804 153694
rect 296204 117694 296804 153458
rect 296204 117458 296386 117694
rect 296622 117458 296804 117694
rect 296204 81694 296804 117458
rect 296204 81458 296386 81694
rect 296622 81458 296804 81694
rect 296204 45694 296804 81458
rect 296204 45458 296386 45694
rect 296622 45458 296804 45694
rect 296204 9694 296804 45458
rect 296204 9458 296386 9694
rect 296622 9458 296804 9694
rect 296204 -4186 296804 9458
rect 296204 -4422 296386 -4186
rect 296622 -4422 296804 -4186
rect 296204 -4506 296804 -4422
rect 296204 -4742 296386 -4506
rect 296622 -4742 296804 -4506
rect 296204 -5734 296804 -4742
rect 299904 697394 300504 710042
rect 317904 711558 318504 711590
rect 317904 711322 318086 711558
rect 318322 711322 318504 711558
rect 317904 711238 318504 711322
rect 317904 711002 318086 711238
rect 318322 711002 318504 711238
rect 314204 709638 314804 709670
rect 314204 709402 314386 709638
rect 314622 709402 314804 709638
rect 314204 709318 314804 709402
rect 314204 709082 314386 709318
rect 314622 709082 314804 709318
rect 310504 707718 311104 707750
rect 310504 707482 310686 707718
rect 310922 707482 311104 707718
rect 310504 707398 311104 707482
rect 310504 707162 310686 707398
rect 310922 707162 311104 707398
rect 299904 697158 300086 697394
rect 300322 697158 300504 697394
rect 299904 661394 300504 697158
rect 299904 661158 300086 661394
rect 300322 661158 300504 661394
rect 299904 625394 300504 661158
rect 299904 625158 300086 625394
rect 300322 625158 300504 625394
rect 299904 589394 300504 625158
rect 299904 589158 300086 589394
rect 300322 589158 300504 589394
rect 299904 553394 300504 589158
rect 299904 553158 300086 553394
rect 300322 553158 300504 553394
rect 299904 517394 300504 553158
rect 299904 517158 300086 517394
rect 300322 517158 300504 517394
rect 299904 481394 300504 517158
rect 299904 481158 300086 481394
rect 300322 481158 300504 481394
rect 299904 445394 300504 481158
rect 299904 445158 300086 445394
rect 300322 445158 300504 445394
rect 299904 409394 300504 445158
rect 299904 409158 300086 409394
rect 300322 409158 300504 409394
rect 299904 373394 300504 409158
rect 299904 373158 300086 373394
rect 300322 373158 300504 373394
rect 299904 337394 300504 373158
rect 299904 337158 300086 337394
rect 300322 337158 300504 337394
rect 299904 301394 300504 337158
rect 299904 301158 300086 301394
rect 300322 301158 300504 301394
rect 299904 265394 300504 301158
rect 299904 265158 300086 265394
rect 300322 265158 300504 265394
rect 299904 229394 300504 265158
rect 299904 229158 300086 229394
rect 300322 229158 300504 229394
rect 299904 193394 300504 229158
rect 299904 193158 300086 193394
rect 300322 193158 300504 193394
rect 299904 157394 300504 193158
rect 299904 157158 300086 157394
rect 300322 157158 300504 157394
rect 299904 121394 300504 157158
rect 299904 121158 300086 121394
rect 300322 121158 300504 121394
rect 299904 85394 300504 121158
rect 299904 85158 300086 85394
rect 300322 85158 300504 85394
rect 299904 49394 300504 85158
rect 299904 49158 300086 49394
rect 300322 49158 300504 49394
rect 299904 13394 300504 49158
rect 299904 13158 300086 13394
rect 300322 13158 300504 13394
rect 281904 -7302 282086 -7066
rect 282322 -7302 282504 -7066
rect 281904 -7386 282504 -7302
rect 281904 -7622 282086 -7386
rect 282322 -7622 282504 -7386
rect 281904 -7654 282504 -7622
rect 299904 -6106 300504 13158
rect 306804 705798 307404 705830
rect 306804 705562 306986 705798
rect 307222 705562 307404 705798
rect 306804 705478 307404 705562
rect 306804 705242 306986 705478
rect 307222 705242 307404 705478
rect 306804 668294 307404 705242
rect 306804 668058 306986 668294
rect 307222 668058 307404 668294
rect 306804 632294 307404 668058
rect 306804 632058 306986 632294
rect 307222 632058 307404 632294
rect 306804 596294 307404 632058
rect 306804 596058 306986 596294
rect 307222 596058 307404 596294
rect 306804 560294 307404 596058
rect 306804 560058 306986 560294
rect 307222 560058 307404 560294
rect 306804 524294 307404 560058
rect 306804 524058 306986 524294
rect 307222 524058 307404 524294
rect 306804 488294 307404 524058
rect 306804 488058 306986 488294
rect 307222 488058 307404 488294
rect 306804 452294 307404 488058
rect 306804 452058 306986 452294
rect 307222 452058 307404 452294
rect 306804 416294 307404 452058
rect 306804 416058 306986 416294
rect 307222 416058 307404 416294
rect 306804 380294 307404 416058
rect 306804 380058 306986 380294
rect 307222 380058 307404 380294
rect 306804 344294 307404 380058
rect 306804 344058 306986 344294
rect 307222 344058 307404 344294
rect 306804 308294 307404 344058
rect 306804 308058 306986 308294
rect 307222 308058 307404 308294
rect 306804 272294 307404 308058
rect 306804 272058 306986 272294
rect 307222 272058 307404 272294
rect 306804 236294 307404 272058
rect 306804 236058 306986 236294
rect 307222 236058 307404 236294
rect 306804 200294 307404 236058
rect 306804 200058 306986 200294
rect 307222 200058 307404 200294
rect 306804 164294 307404 200058
rect 306804 164058 306986 164294
rect 307222 164058 307404 164294
rect 306804 128294 307404 164058
rect 306804 128058 306986 128294
rect 307222 128058 307404 128294
rect 306804 92294 307404 128058
rect 306804 92058 306986 92294
rect 307222 92058 307404 92294
rect 306804 56294 307404 92058
rect 306804 56058 306986 56294
rect 307222 56058 307404 56294
rect 306804 20294 307404 56058
rect 306804 20058 306986 20294
rect 307222 20058 307404 20294
rect 306804 -1306 307404 20058
rect 306804 -1542 306986 -1306
rect 307222 -1542 307404 -1306
rect 306804 -1626 307404 -1542
rect 306804 -1862 306986 -1626
rect 307222 -1862 307404 -1626
rect 306804 -1894 307404 -1862
rect 310504 671994 311104 707162
rect 310504 671758 310686 671994
rect 310922 671758 311104 671994
rect 310504 635994 311104 671758
rect 310504 635758 310686 635994
rect 310922 635758 311104 635994
rect 310504 599994 311104 635758
rect 310504 599758 310686 599994
rect 310922 599758 311104 599994
rect 310504 563994 311104 599758
rect 310504 563758 310686 563994
rect 310922 563758 311104 563994
rect 310504 527994 311104 563758
rect 310504 527758 310686 527994
rect 310922 527758 311104 527994
rect 310504 491994 311104 527758
rect 310504 491758 310686 491994
rect 310922 491758 311104 491994
rect 310504 455994 311104 491758
rect 310504 455758 310686 455994
rect 310922 455758 311104 455994
rect 310504 419994 311104 455758
rect 310504 419758 310686 419994
rect 310922 419758 311104 419994
rect 310504 383994 311104 419758
rect 310504 383758 310686 383994
rect 310922 383758 311104 383994
rect 310504 347994 311104 383758
rect 310504 347758 310686 347994
rect 310922 347758 311104 347994
rect 310504 311994 311104 347758
rect 310504 311758 310686 311994
rect 310922 311758 311104 311994
rect 310504 275994 311104 311758
rect 310504 275758 310686 275994
rect 310922 275758 311104 275994
rect 310504 239994 311104 275758
rect 310504 239758 310686 239994
rect 310922 239758 311104 239994
rect 310504 203994 311104 239758
rect 310504 203758 310686 203994
rect 310922 203758 311104 203994
rect 310504 167994 311104 203758
rect 310504 167758 310686 167994
rect 310922 167758 311104 167994
rect 310504 131994 311104 167758
rect 310504 131758 310686 131994
rect 310922 131758 311104 131994
rect 310504 95994 311104 131758
rect 310504 95758 310686 95994
rect 310922 95758 311104 95994
rect 310504 59994 311104 95758
rect 310504 59758 310686 59994
rect 310922 59758 311104 59994
rect 310504 23994 311104 59758
rect 310504 23758 310686 23994
rect 310922 23758 311104 23994
rect 310504 -3226 311104 23758
rect 310504 -3462 310686 -3226
rect 310922 -3462 311104 -3226
rect 310504 -3546 311104 -3462
rect 310504 -3782 310686 -3546
rect 310922 -3782 311104 -3546
rect 310504 -3814 311104 -3782
rect 314204 675694 314804 709082
rect 314204 675458 314386 675694
rect 314622 675458 314804 675694
rect 314204 639694 314804 675458
rect 314204 639458 314386 639694
rect 314622 639458 314804 639694
rect 314204 603694 314804 639458
rect 314204 603458 314386 603694
rect 314622 603458 314804 603694
rect 314204 567694 314804 603458
rect 314204 567458 314386 567694
rect 314622 567458 314804 567694
rect 314204 531694 314804 567458
rect 314204 531458 314386 531694
rect 314622 531458 314804 531694
rect 314204 495694 314804 531458
rect 314204 495458 314386 495694
rect 314622 495458 314804 495694
rect 314204 459694 314804 495458
rect 314204 459458 314386 459694
rect 314622 459458 314804 459694
rect 314204 423694 314804 459458
rect 314204 423458 314386 423694
rect 314622 423458 314804 423694
rect 314204 387694 314804 423458
rect 314204 387458 314386 387694
rect 314622 387458 314804 387694
rect 314204 351694 314804 387458
rect 314204 351458 314386 351694
rect 314622 351458 314804 351694
rect 314204 315694 314804 351458
rect 314204 315458 314386 315694
rect 314622 315458 314804 315694
rect 314204 279694 314804 315458
rect 314204 279458 314386 279694
rect 314622 279458 314804 279694
rect 314204 243694 314804 279458
rect 314204 243458 314386 243694
rect 314622 243458 314804 243694
rect 314204 207694 314804 243458
rect 314204 207458 314386 207694
rect 314622 207458 314804 207694
rect 314204 171694 314804 207458
rect 314204 171458 314386 171694
rect 314622 171458 314804 171694
rect 314204 135694 314804 171458
rect 314204 135458 314386 135694
rect 314622 135458 314804 135694
rect 314204 99694 314804 135458
rect 314204 99458 314386 99694
rect 314622 99458 314804 99694
rect 314204 63694 314804 99458
rect 314204 63458 314386 63694
rect 314622 63458 314804 63694
rect 314204 27694 314804 63458
rect 314204 27458 314386 27694
rect 314622 27458 314804 27694
rect 314204 -5146 314804 27458
rect 314204 -5382 314386 -5146
rect 314622 -5382 314804 -5146
rect 314204 -5466 314804 -5382
rect 314204 -5702 314386 -5466
rect 314622 -5702 314804 -5466
rect 314204 -5734 314804 -5702
rect 317904 679394 318504 711002
rect 335904 710598 336504 711590
rect 335904 710362 336086 710598
rect 336322 710362 336504 710598
rect 335904 710278 336504 710362
rect 335904 710042 336086 710278
rect 336322 710042 336504 710278
rect 332204 708678 332804 709670
rect 332204 708442 332386 708678
rect 332622 708442 332804 708678
rect 332204 708358 332804 708442
rect 332204 708122 332386 708358
rect 332622 708122 332804 708358
rect 328504 706758 329104 707750
rect 328504 706522 328686 706758
rect 328922 706522 329104 706758
rect 328504 706438 329104 706522
rect 328504 706202 328686 706438
rect 328922 706202 329104 706438
rect 317904 679158 318086 679394
rect 318322 679158 318504 679394
rect 317904 643394 318504 679158
rect 317904 643158 318086 643394
rect 318322 643158 318504 643394
rect 317904 607394 318504 643158
rect 317904 607158 318086 607394
rect 318322 607158 318504 607394
rect 317904 571394 318504 607158
rect 317904 571158 318086 571394
rect 318322 571158 318504 571394
rect 317904 535394 318504 571158
rect 317904 535158 318086 535394
rect 318322 535158 318504 535394
rect 317904 499394 318504 535158
rect 317904 499158 318086 499394
rect 318322 499158 318504 499394
rect 317904 463394 318504 499158
rect 317904 463158 318086 463394
rect 318322 463158 318504 463394
rect 317904 427394 318504 463158
rect 317904 427158 318086 427394
rect 318322 427158 318504 427394
rect 317904 391394 318504 427158
rect 317904 391158 318086 391394
rect 318322 391158 318504 391394
rect 317904 355394 318504 391158
rect 317904 355158 318086 355394
rect 318322 355158 318504 355394
rect 317904 319394 318504 355158
rect 317904 319158 318086 319394
rect 318322 319158 318504 319394
rect 317904 283394 318504 319158
rect 317904 283158 318086 283394
rect 318322 283158 318504 283394
rect 317904 247394 318504 283158
rect 317904 247158 318086 247394
rect 318322 247158 318504 247394
rect 317904 211394 318504 247158
rect 317904 211158 318086 211394
rect 318322 211158 318504 211394
rect 317904 175394 318504 211158
rect 317904 175158 318086 175394
rect 318322 175158 318504 175394
rect 317904 139394 318504 175158
rect 317904 139158 318086 139394
rect 318322 139158 318504 139394
rect 317904 103394 318504 139158
rect 317904 103158 318086 103394
rect 318322 103158 318504 103394
rect 317904 67394 318504 103158
rect 317904 67158 318086 67394
rect 318322 67158 318504 67394
rect 317904 31394 318504 67158
rect 317904 31158 318086 31394
rect 318322 31158 318504 31394
rect 299904 -6342 300086 -6106
rect 300322 -6342 300504 -6106
rect 299904 -6426 300504 -6342
rect 299904 -6662 300086 -6426
rect 300322 -6662 300504 -6426
rect 299904 -7654 300504 -6662
rect 317904 -7066 318504 31158
rect 324804 704838 325404 705830
rect 324804 704602 324986 704838
rect 325222 704602 325404 704838
rect 324804 704518 325404 704602
rect 324804 704282 324986 704518
rect 325222 704282 325404 704518
rect 324804 686294 325404 704282
rect 324804 686058 324986 686294
rect 325222 686058 325404 686294
rect 324804 650294 325404 686058
rect 324804 650058 324986 650294
rect 325222 650058 325404 650294
rect 324804 614294 325404 650058
rect 324804 614058 324986 614294
rect 325222 614058 325404 614294
rect 324804 578294 325404 614058
rect 324804 578058 324986 578294
rect 325222 578058 325404 578294
rect 324804 542294 325404 578058
rect 324804 542058 324986 542294
rect 325222 542058 325404 542294
rect 324804 506294 325404 542058
rect 324804 506058 324986 506294
rect 325222 506058 325404 506294
rect 324804 470294 325404 506058
rect 324804 470058 324986 470294
rect 325222 470058 325404 470294
rect 324804 434294 325404 470058
rect 324804 434058 324986 434294
rect 325222 434058 325404 434294
rect 324804 398294 325404 434058
rect 324804 398058 324986 398294
rect 325222 398058 325404 398294
rect 324804 362294 325404 398058
rect 324804 362058 324986 362294
rect 325222 362058 325404 362294
rect 324804 326294 325404 362058
rect 324804 326058 324986 326294
rect 325222 326058 325404 326294
rect 324804 290294 325404 326058
rect 324804 290058 324986 290294
rect 325222 290058 325404 290294
rect 324804 254294 325404 290058
rect 324804 254058 324986 254294
rect 325222 254058 325404 254294
rect 324804 218294 325404 254058
rect 324804 218058 324986 218294
rect 325222 218058 325404 218294
rect 324804 182294 325404 218058
rect 324804 182058 324986 182294
rect 325222 182058 325404 182294
rect 324804 146294 325404 182058
rect 324804 146058 324986 146294
rect 325222 146058 325404 146294
rect 324804 110294 325404 146058
rect 324804 110058 324986 110294
rect 325222 110058 325404 110294
rect 324804 74294 325404 110058
rect 324804 74058 324986 74294
rect 325222 74058 325404 74294
rect 324804 38294 325404 74058
rect 324804 38058 324986 38294
rect 325222 38058 325404 38294
rect 324804 2294 325404 38058
rect 324804 2058 324986 2294
rect 325222 2058 325404 2294
rect 324804 -346 325404 2058
rect 324804 -582 324986 -346
rect 325222 -582 325404 -346
rect 324804 -666 325404 -582
rect 324804 -902 324986 -666
rect 325222 -902 325404 -666
rect 324804 -1894 325404 -902
rect 328504 689994 329104 706202
rect 328504 689758 328686 689994
rect 328922 689758 329104 689994
rect 328504 653994 329104 689758
rect 328504 653758 328686 653994
rect 328922 653758 329104 653994
rect 328504 617994 329104 653758
rect 328504 617758 328686 617994
rect 328922 617758 329104 617994
rect 328504 581994 329104 617758
rect 328504 581758 328686 581994
rect 328922 581758 329104 581994
rect 328504 545994 329104 581758
rect 328504 545758 328686 545994
rect 328922 545758 329104 545994
rect 328504 509994 329104 545758
rect 328504 509758 328686 509994
rect 328922 509758 329104 509994
rect 328504 473994 329104 509758
rect 328504 473758 328686 473994
rect 328922 473758 329104 473994
rect 328504 437994 329104 473758
rect 328504 437758 328686 437994
rect 328922 437758 329104 437994
rect 328504 401994 329104 437758
rect 328504 401758 328686 401994
rect 328922 401758 329104 401994
rect 328504 365994 329104 401758
rect 328504 365758 328686 365994
rect 328922 365758 329104 365994
rect 328504 329994 329104 365758
rect 328504 329758 328686 329994
rect 328922 329758 329104 329994
rect 328504 293994 329104 329758
rect 328504 293758 328686 293994
rect 328922 293758 329104 293994
rect 328504 257994 329104 293758
rect 328504 257758 328686 257994
rect 328922 257758 329104 257994
rect 328504 221994 329104 257758
rect 328504 221758 328686 221994
rect 328922 221758 329104 221994
rect 328504 185994 329104 221758
rect 328504 185758 328686 185994
rect 328922 185758 329104 185994
rect 328504 149994 329104 185758
rect 328504 149758 328686 149994
rect 328922 149758 329104 149994
rect 328504 113994 329104 149758
rect 328504 113758 328686 113994
rect 328922 113758 329104 113994
rect 328504 77994 329104 113758
rect 328504 77758 328686 77994
rect 328922 77758 329104 77994
rect 328504 41994 329104 77758
rect 328504 41758 328686 41994
rect 328922 41758 329104 41994
rect 328504 5994 329104 41758
rect 328504 5758 328686 5994
rect 328922 5758 329104 5994
rect 328504 -2266 329104 5758
rect 328504 -2502 328686 -2266
rect 328922 -2502 329104 -2266
rect 328504 -2586 329104 -2502
rect 328504 -2822 328686 -2586
rect 328922 -2822 329104 -2586
rect 328504 -3814 329104 -2822
rect 332204 693694 332804 708122
rect 332204 693458 332386 693694
rect 332622 693458 332804 693694
rect 332204 657694 332804 693458
rect 332204 657458 332386 657694
rect 332622 657458 332804 657694
rect 332204 621694 332804 657458
rect 332204 621458 332386 621694
rect 332622 621458 332804 621694
rect 332204 585694 332804 621458
rect 332204 585458 332386 585694
rect 332622 585458 332804 585694
rect 332204 549694 332804 585458
rect 332204 549458 332386 549694
rect 332622 549458 332804 549694
rect 332204 513694 332804 549458
rect 332204 513458 332386 513694
rect 332622 513458 332804 513694
rect 332204 477694 332804 513458
rect 332204 477458 332386 477694
rect 332622 477458 332804 477694
rect 332204 441694 332804 477458
rect 332204 441458 332386 441694
rect 332622 441458 332804 441694
rect 332204 405694 332804 441458
rect 332204 405458 332386 405694
rect 332622 405458 332804 405694
rect 332204 369694 332804 405458
rect 332204 369458 332386 369694
rect 332622 369458 332804 369694
rect 332204 333694 332804 369458
rect 332204 333458 332386 333694
rect 332622 333458 332804 333694
rect 332204 297694 332804 333458
rect 332204 297458 332386 297694
rect 332622 297458 332804 297694
rect 332204 261694 332804 297458
rect 332204 261458 332386 261694
rect 332622 261458 332804 261694
rect 332204 225694 332804 261458
rect 332204 225458 332386 225694
rect 332622 225458 332804 225694
rect 332204 189694 332804 225458
rect 332204 189458 332386 189694
rect 332622 189458 332804 189694
rect 332204 153694 332804 189458
rect 332204 153458 332386 153694
rect 332622 153458 332804 153694
rect 332204 117694 332804 153458
rect 332204 117458 332386 117694
rect 332622 117458 332804 117694
rect 332204 81694 332804 117458
rect 332204 81458 332386 81694
rect 332622 81458 332804 81694
rect 332204 45694 332804 81458
rect 332204 45458 332386 45694
rect 332622 45458 332804 45694
rect 332204 9694 332804 45458
rect 332204 9458 332386 9694
rect 332622 9458 332804 9694
rect 332204 -4186 332804 9458
rect 332204 -4422 332386 -4186
rect 332622 -4422 332804 -4186
rect 332204 -4506 332804 -4422
rect 332204 -4742 332386 -4506
rect 332622 -4742 332804 -4506
rect 332204 -5734 332804 -4742
rect 335904 697394 336504 710042
rect 353904 711558 354504 711590
rect 353904 711322 354086 711558
rect 354322 711322 354504 711558
rect 353904 711238 354504 711322
rect 353904 711002 354086 711238
rect 354322 711002 354504 711238
rect 350204 709638 350804 709670
rect 350204 709402 350386 709638
rect 350622 709402 350804 709638
rect 350204 709318 350804 709402
rect 350204 709082 350386 709318
rect 350622 709082 350804 709318
rect 346504 707718 347104 707750
rect 346504 707482 346686 707718
rect 346922 707482 347104 707718
rect 346504 707398 347104 707482
rect 346504 707162 346686 707398
rect 346922 707162 347104 707398
rect 335904 697158 336086 697394
rect 336322 697158 336504 697394
rect 335904 661394 336504 697158
rect 335904 661158 336086 661394
rect 336322 661158 336504 661394
rect 335904 625394 336504 661158
rect 335904 625158 336086 625394
rect 336322 625158 336504 625394
rect 335904 589394 336504 625158
rect 335904 589158 336086 589394
rect 336322 589158 336504 589394
rect 335904 553394 336504 589158
rect 335904 553158 336086 553394
rect 336322 553158 336504 553394
rect 335904 517394 336504 553158
rect 335904 517158 336086 517394
rect 336322 517158 336504 517394
rect 335904 481394 336504 517158
rect 335904 481158 336086 481394
rect 336322 481158 336504 481394
rect 335904 445394 336504 481158
rect 335904 445158 336086 445394
rect 336322 445158 336504 445394
rect 335904 409394 336504 445158
rect 342804 705798 343404 705830
rect 342804 705562 342986 705798
rect 343222 705562 343404 705798
rect 342804 705478 343404 705562
rect 342804 705242 342986 705478
rect 343222 705242 343404 705478
rect 342804 668294 343404 705242
rect 342804 668058 342986 668294
rect 343222 668058 343404 668294
rect 342804 632294 343404 668058
rect 342804 632058 342986 632294
rect 343222 632058 343404 632294
rect 342804 596294 343404 632058
rect 342804 596058 342986 596294
rect 343222 596058 343404 596294
rect 342804 560294 343404 596058
rect 342804 560058 342986 560294
rect 343222 560058 343404 560294
rect 342804 524294 343404 560058
rect 342804 524058 342986 524294
rect 343222 524058 343404 524294
rect 342804 488294 343404 524058
rect 342804 488058 342986 488294
rect 343222 488058 343404 488294
rect 342804 452294 343404 488058
rect 342804 452058 342986 452294
rect 343222 452058 343404 452294
rect 342804 425308 343404 452058
rect 346504 671994 347104 707162
rect 346504 671758 346686 671994
rect 346922 671758 347104 671994
rect 346504 635994 347104 671758
rect 346504 635758 346686 635994
rect 346922 635758 347104 635994
rect 346504 599994 347104 635758
rect 346504 599758 346686 599994
rect 346922 599758 347104 599994
rect 346504 563994 347104 599758
rect 346504 563758 346686 563994
rect 346922 563758 347104 563994
rect 346504 527994 347104 563758
rect 346504 527758 346686 527994
rect 346922 527758 347104 527994
rect 346504 491994 347104 527758
rect 346504 491758 346686 491994
rect 346922 491758 347104 491994
rect 346504 455994 347104 491758
rect 346504 455758 346686 455994
rect 346922 455758 347104 455994
rect 346504 425308 347104 455758
rect 350204 675694 350804 709082
rect 350204 675458 350386 675694
rect 350622 675458 350804 675694
rect 350204 639694 350804 675458
rect 350204 639458 350386 639694
rect 350622 639458 350804 639694
rect 350204 603694 350804 639458
rect 350204 603458 350386 603694
rect 350622 603458 350804 603694
rect 350204 567694 350804 603458
rect 350204 567458 350386 567694
rect 350622 567458 350804 567694
rect 350204 531694 350804 567458
rect 350204 531458 350386 531694
rect 350622 531458 350804 531694
rect 350204 495694 350804 531458
rect 350204 495458 350386 495694
rect 350622 495458 350804 495694
rect 350204 459694 350804 495458
rect 350204 459458 350386 459694
rect 350622 459458 350804 459694
rect 350204 425308 350804 459458
rect 353904 679394 354504 711002
rect 371904 710598 372504 711590
rect 371904 710362 372086 710598
rect 372322 710362 372504 710598
rect 371904 710278 372504 710362
rect 371904 710042 372086 710278
rect 372322 710042 372504 710278
rect 368204 708678 368804 709670
rect 368204 708442 368386 708678
rect 368622 708442 368804 708678
rect 368204 708358 368804 708442
rect 368204 708122 368386 708358
rect 368622 708122 368804 708358
rect 364504 706758 365104 707750
rect 364504 706522 364686 706758
rect 364922 706522 365104 706758
rect 364504 706438 365104 706522
rect 364504 706202 364686 706438
rect 364922 706202 365104 706438
rect 353904 679158 354086 679394
rect 354322 679158 354504 679394
rect 353904 643394 354504 679158
rect 353904 643158 354086 643394
rect 354322 643158 354504 643394
rect 353904 607394 354504 643158
rect 353904 607158 354086 607394
rect 354322 607158 354504 607394
rect 353904 571394 354504 607158
rect 353904 571158 354086 571394
rect 354322 571158 354504 571394
rect 353904 535394 354504 571158
rect 353904 535158 354086 535394
rect 354322 535158 354504 535394
rect 353904 499394 354504 535158
rect 353904 499158 354086 499394
rect 354322 499158 354504 499394
rect 353904 463394 354504 499158
rect 353904 463158 354086 463394
rect 354322 463158 354504 463394
rect 353904 427394 354504 463158
rect 353904 427158 354086 427394
rect 354322 427158 354504 427394
rect 353904 425308 354504 427158
rect 360804 704838 361404 705830
rect 360804 704602 360986 704838
rect 361222 704602 361404 704838
rect 360804 704518 361404 704602
rect 360804 704282 360986 704518
rect 361222 704282 361404 704518
rect 360804 686294 361404 704282
rect 360804 686058 360986 686294
rect 361222 686058 361404 686294
rect 360804 650294 361404 686058
rect 360804 650058 360986 650294
rect 361222 650058 361404 650294
rect 360804 614294 361404 650058
rect 360804 614058 360986 614294
rect 361222 614058 361404 614294
rect 360804 578294 361404 614058
rect 360804 578058 360986 578294
rect 361222 578058 361404 578294
rect 360804 542294 361404 578058
rect 360804 542058 360986 542294
rect 361222 542058 361404 542294
rect 360804 506294 361404 542058
rect 360804 506058 360986 506294
rect 361222 506058 361404 506294
rect 360804 470294 361404 506058
rect 360804 470058 360986 470294
rect 361222 470058 361404 470294
rect 360804 434294 361404 470058
rect 360804 434058 360986 434294
rect 361222 434058 361404 434294
rect 360804 425308 361404 434058
rect 364504 689994 365104 706202
rect 364504 689758 364686 689994
rect 364922 689758 365104 689994
rect 364504 653994 365104 689758
rect 364504 653758 364686 653994
rect 364922 653758 365104 653994
rect 364504 617994 365104 653758
rect 364504 617758 364686 617994
rect 364922 617758 365104 617994
rect 364504 581994 365104 617758
rect 364504 581758 364686 581994
rect 364922 581758 365104 581994
rect 364504 545994 365104 581758
rect 364504 545758 364686 545994
rect 364922 545758 365104 545994
rect 364504 509994 365104 545758
rect 364504 509758 364686 509994
rect 364922 509758 365104 509994
rect 364504 473994 365104 509758
rect 364504 473758 364686 473994
rect 364922 473758 365104 473994
rect 364504 437994 365104 473758
rect 364504 437758 364686 437994
rect 364922 437758 365104 437994
rect 364504 425308 365104 437758
rect 368204 693694 368804 708122
rect 368204 693458 368386 693694
rect 368622 693458 368804 693694
rect 368204 657694 368804 693458
rect 368204 657458 368386 657694
rect 368622 657458 368804 657694
rect 368204 621694 368804 657458
rect 368204 621458 368386 621694
rect 368622 621458 368804 621694
rect 368204 585694 368804 621458
rect 368204 585458 368386 585694
rect 368622 585458 368804 585694
rect 368204 549694 368804 585458
rect 368204 549458 368386 549694
rect 368622 549458 368804 549694
rect 368204 513694 368804 549458
rect 368204 513458 368386 513694
rect 368622 513458 368804 513694
rect 368204 477694 368804 513458
rect 368204 477458 368386 477694
rect 368622 477458 368804 477694
rect 368204 441694 368804 477458
rect 368204 441458 368386 441694
rect 368622 441458 368804 441694
rect 368204 425308 368804 441458
rect 371904 697394 372504 710042
rect 389904 711558 390504 711590
rect 389904 711322 390086 711558
rect 390322 711322 390504 711558
rect 389904 711238 390504 711322
rect 389904 711002 390086 711238
rect 390322 711002 390504 711238
rect 386204 709638 386804 709670
rect 386204 709402 386386 709638
rect 386622 709402 386804 709638
rect 386204 709318 386804 709402
rect 386204 709082 386386 709318
rect 386622 709082 386804 709318
rect 382504 707718 383104 707750
rect 382504 707482 382686 707718
rect 382922 707482 383104 707718
rect 382504 707398 383104 707482
rect 382504 707162 382686 707398
rect 382922 707162 383104 707398
rect 371904 697158 372086 697394
rect 372322 697158 372504 697394
rect 371904 661394 372504 697158
rect 371904 661158 372086 661394
rect 372322 661158 372504 661394
rect 371904 625394 372504 661158
rect 371904 625158 372086 625394
rect 372322 625158 372504 625394
rect 371904 589394 372504 625158
rect 371904 589158 372086 589394
rect 372322 589158 372504 589394
rect 371904 553394 372504 589158
rect 371904 553158 372086 553394
rect 372322 553158 372504 553394
rect 371904 517394 372504 553158
rect 371904 517158 372086 517394
rect 372322 517158 372504 517394
rect 371904 481394 372504 517158
rect 371904 481158 372086 481394
rect 372322 481158 372504 481394
rect 371904 445394 372504 481158
rect 371904 445158 372086 445394
rect 372322 445158 372504 445394
rect 371904 425308 372504 445158
rect 378804 705798 379404 705830
rect 378804 705562 378986 705798
rect 379222 705562 379404 705798
rect 378804 705478 379404 705562
rect 378804 705242 378986 705478
rect 379222 705242 379404 705478
rect 378804 668294 379404 705242
rect 378804 668058 378986 668294
rect 379222 668058 379404 668294
rect 378804 632294 379404 668058
rect 378804 632058 378986 632294
rect 379222 632058 379404 632294
rect 378804 596294 379404 632058
rect 378804 596058 378986 596294
rect 379222 596058 379404 596294
rect 378804 560294 379404 596058
rect 378804 560058 378986 560294
rect 379222 560058 379404 560294
rect 378804 524294 379404 560058
rect 378804 524058 378986 524294
rect 379222 524058 379404 524294
rect 378804 488294 379404 524058
rect 378804 488058 378986 488294
rect 379222 488058 379404 488294
rect 378804 452294 379404 488058
rect 378804 452058 378986 452294
rect 379222 452058 379404 452294
rect 378804 425308 379404 452058
rect 382504 671994 383104 707162
rect 382504 671758 382686 671994
rect 382922 671758 383104 671994
rect 382504 635994 383104 671758
rect 382504 635758 382686 635994
rect 382922 635758 383104 635994
rect 382504 599994 383104 635758
rect 382504 599758 382686 599994
rect 382922 599758 383104 599994
rect 382504 563994 383104 599758
rect 382504 563758 382686 563994
rect 382922 563758 383104 563994
rect 382504 527994 383104 563758
rect 382504 527758 382686 527994
rect 382922 527758 383104 527994
rect 382504 491994 383104 527758
rect 382504 491758 382686 491994
rect 382922 491758 383104 491994
rect 382504 455994 383104 491758
rect 382504 455758 382686 455994
rect 382922 455758 383104 455994
rect 382504 425308 383104 455758
rect 386204 675694 386804 709082
rect 386204 675458 386386 675694
rect 386622 675458 386804 675694
rect 386204 639694 386804 675458
rect 386204 639458 386386 639694
rect 386622 639458 386804 639694
rect 386204 603694 386804 639458
rect 386204 603458 386386 603694
rect 386622 603458 386804 603694
rect 386204 567694 386804 603458
rect 386204 567458 386386 567694
rect 386622 567458 386804 567694
rect 386204 531694 386804 567458
rect 386204 531458 386386 531694
rect 386622 531458 386804 531694
rect 386204 495694 386804 531458
rect 386204 495458 386386 495694
rect 386622 495458 386804 495694
rect 386204 459694 386804 495458
rect 386204 459458 386386 459694
rect 386622 459458 386804 459694
rect 386204 425308 386804 459458
rect 389904 679394 390504 711002
rect 407904 710598 408504 711590
rect 407904 710362 408086 710598
rect 408322 710362 408504 710598
rect 407904 710278 408504 710362
rect 407904 710042 408086 710278
rect 408322 710042 408504 710278
rect 404204 708678 404804 709670
rect 404204 708442 404386 708678
rect 404622 708442 404804 708678
rect 404204 708358 404804 708442
rect 404204 708122 404386 708358
rect 404622 708122 404804 708358
rect 400504 706758 401104 707750
rect 400504 706522 400686 706758
rect 400922 706522 401104 706758
rect 400504 706438 401104 706522
rect 400504 706202 400686 706438
rect 400922 706202 401104 706438
rect 389904 679158 390086 679394
rect 390322 679158 390504 679394
rect 389904 643394 390504 679158
rect 389904 643158 390086 643394
rect 390322 643158 390504 643394
rect 389904 607394 390504 643158
rect 389904 607158 390086 607394
rect 390322 607158 390504 607394
rect 389904 571394 390504 607158
rect 389904 571158 390086 571394
rect 390322 571158 390504 571394
rect 389904 535394 390504 571158
rect 389904 535158 390086 535394
rect 390322 535158 390504 535394
rect 389904 499394 390504 535158
rect 389904 499158 390086 499394
rect 390322 499158 390504 499394
rect 389904 463394 390504 499158
rect 389904 463158 390086 463394
rect 390322 463158 390504 463394
rect 389904 427394 390504 463158
rect 389904 427158 390086 427394
rect 390322 427158 390504 427394
rect 389904 425308 390504 427158
rect 396804 704838 397404 705830
rect 396804 704602 396986 704838
rect 397222 704602 397404 704838
rect 396804 704518 397404 704602
rect 396804 704282 396986 704518
rect 397222 704282 397404 704518
rect 396804 686294 397404 704282
rect 396804 686058 396986 686294
rect 397222 686058 397404 686294
rect 396804 650294 397404 686058
rect 396804 650058 396986 650294
rect 397222 650058 397404 650294
rect 396804 614294 397404 650058
rect 396804 614058 396986 614294
rect 397222 614058 397404 614294
rect 396804 578294 397404 614058
rect 396804 578058 396986 578294
rect 397222 578058 397404 578294
rect 396804 542294 397404 578058
rect 396804 542058 396986 542294
rect 397222 542058 397404 542294
rect 396804 506294 397404 542058
rect 396804 506058 396986 506294
rect 397222 506058 397404 506294
rect 396804 470294 397404 506058
rect 396804 470058 396986 470294
rect 397222 470058 397404 470294
rect 396804 434294 397404 470058
rect 396804 434058 396986 434294
rect 397222 434058 397404 434294
rect 396804 425308 397404 434058
rect 400504 689994 401104 706202
rect 400504 689758 400686 689994
rect 400922 689758 401104 689994
rect 400504 653994 401104 689758
rect 400504 653758 400686 653994
rect 400922 653758 401104 653994
rect 400504 617994 401104 653758
rect 400504 617758 400686 617994
rect 400922 617758 401104 617994
rect 400504 581994 401104 617758
rect 400504 581758 400686 581994
rect 400922 581758 401104 581994
rect 400504 545994 401104 581758
rect 400504 545758 400686 545994
rect 400922 545758 401104 545994
rect 400504 509994 401104 545758
rect 400504 509758 400686 509994
rect 400922 509758 401104 509994
rect 400504 473994 401104 509758
rect 400504 473758 400686 473994
rect 400922 473758 401104 473994
rect 400504 437994 401104 473758
rect 400504 437758 400686 437994
rect 400922 437758 401104 437994
rect 400504 425308 401104 437758
rect 404204 693694 404804 708122
rect 404204 693458 404386 693694
rect 404622 693458 404804 693694
rect 404204 657694 404804 693458
rect 404204 657458 404386 657694
rect 404622 657458 404804 657694
rect 404204 621694 404804 657458
rect 404204 621458 404386 621694
rect 404622 621458 404804 621694
rect 404204 585694 404804 621458
rect 404204 585458 404386 585694
rect 404622 585458 404804 585694
rect 404204 549694 404804 585458
rect 404204 549458 404386 549694
rect 404622 549458 404804 549694
rect 404204 513694 404804 549458
rect 404204 513458 404386 513694
rect 404622 513458 404804 513694
rect 404204 477694 404804 513458
rect 404204 477458 404386 477694
rect 404622 477458 404804 477694
rect 404204 441694 404804 477458
rect 404204 441458 404386 441694
rect 404622 441458 404804 441694
rect 404204 425308 404804 441458
rect 407904 697394 408504 710042
rect 425904 711558 426504 711590
rect 425904 711322 426086 711558
rect 426322 711322 426504 711558
rect 425904 711238 426504 711322
rect 425904 711002 426086 711238
rect 426322 711002 426504 711238
rect 422204 709638 422804 709670
rect 422204 709402 422386 709638
rect 422622 709402 422804 709638
rect 422204 709318 422804 709402
rect 422204 709082 422386 709318
rect 422622 709082 422804 709318
rect 418504 707718 419104 707750
rect 418504 707482 418686 707718
rect 418922 707482 419104 707718
rect 418504 707398 419104 707482
rect 418504 707162 418686 707398
rect 418922 707162 419104 707398
rect 407904 697158 408086 697394
rect 408322 697158 408504 697394
rect 407904 661394 408504 697158
rect 407904 661158 408086 661394
rect 408322 661158 408504 661394
rect 407904 625394 408504 661158
rect 407904 625158 408086 625394
rect 408322 625158 408504 625394
rect 407904 589394 408504 625158
rect 407904 589158 408086 589394
rect 408322 589158 408504 589394
rect 407904 553394 408504 589158
rect 407904 553158 408086 553394
rect 408322 553158 408504 553394
rect 407904 517394 408504 553158
rect 407904 517158 408086 517394
rect 408322 517158 408504 517394
rect 407904 481394 408504 517158
rect 407904 481158 408086 481394
rect 408322 481158 408504 481394
rect 407904 445394 408504 481158
rect 407904 445158 408086 445394
rect 408322 445158 408504 445394
rect 407904 425308 408504 445158
rect 414804 705798 415404 705830
rect 414804 705562 414986 705798
rect 415222 705562 415404 705798
rect 414804 705478 415404 705562
rect 414804 705242 414986 705478
rect 415222 705242 415404 705478
rect 414804 668294 415404 705242
rect 414804 668058 414986 668294
rect 415222 668058 415404 668294
rect 414804 632294 415404 668058
rect 414804 632058 414986 632294
rect 415222 632058 415404 632294
rect 414804 596294 415404 632058
rect 414804 596058 414986 596294
rect 415222 596058 415404 596294
rect 414804 560294 415404 596058
rect 414804 560058 414986 560294
rect 415222 560058 415404 560294
rect 414804 524294 415404 560058
rect 414804 524058 414986 524294
rect 415222 524058 415404 524294
rect 414804 488294 415404 524058
rect 414804 488058 414986 488294
rect 415222 488058 415404 488294
rect 414804 452294 415404 488058
rect 414804 452058 414986 452294
rect 415222 452058 415404 452294
rect 414804 425308 415404 452058
rect 418504 671994 419104 707162
rect 418504 671758 418686 671994
rect 418922 671758 419104 671994
rect 418504 635994 419104 671758
rect 418504 635758 418686 635994
rect 418922 635758 419104 635994
rect 418504 599994 419104 635758
rect 418504 599758 418686 599994
rect 418922 599758 419104 599994
rect 418504 563994 419104 599758
rect 418504 563758 418686 563994
rect 418922 563758 419104 563994
rect 418504 527994 419104 563758
rect 418504 527758 418686 527994
rect 418922 527758 419104 527994
rect 418504 491994 419104 527758
rect 418504 491758 418686 491994
rect 418922 491758 419104 491994
rect 418504 455994 419104 491758
rect 418504 455758 418686 455994
rect 418922 455758 419104 455994
rect 418504 425308 419104 455758
rect 422204 675694 422804 709082
rect 422204 675458 422386 675694
rect 422622 675458 422804 675694
rect 422204 639694 422804 675458
rect 422204 639458 422386 639694
rect 422622 639458 422804 639694
rect 422204 603694 422804 639458
rect 422204 603458 422386 603694
rect 422622 603458 422804 603694
rect 422204 567694 422804 603458
rect 422204 567458 422386 567694
rect 422622 567458 422804 567694
rect 422204 531694 422804 567458
rect 422204 531458 422386 531694
rect 422622 531458 422804 531694
rect 422204 495694 422804 531458
rect 422204 495458 422386 495694
rect 422622 495458 422804 495694
rect 422204 459694 422804 495458
rect 422204 459458 422386 459694
rect 422622 459458 422804 459694
rect 422204 425308 422804 459458
rect 425904 679394 426504 711002
rect 443904 710598 444504 711590
rect 443904 710362 444086 710598
rect 444322 710362 444504 710598
rect 443904 710278 444504 710362
rect 443904 710042 444086 710278
rect 444322 710042 444504 710278
rect 440204 708678 440804 709670
rect 440204 708442 440386 708678
rect 440622 708442 440804 708678
rect 440204 708358 440804 708442
rect 440204 708122 440386 708358
rect 440622 708122 440804 708358
rect 436504 706758 437104 707750
rect 436504 706522 436686 706758
rect 436922 706522 437104 706758
rect 436504 706438 437104 706522
rect 436504 706202 436686 706438
rect 436922 706202 437104 706438
rect 425904 679158 426086 679394
rect 426322 679158 426504 679394
rect 425904 643394 426504 679158
rect 425904 643158 426086 643394
rect 426322 643158 426504 643394
rect 425904 607394 426504 643158
rect 425904 607158 426086 607394
rect 426322 607158 426504 607394
rect 425904 571394 426504 607158
rect 425904 571158 426086 571394
rect 426322 571158 426504 571394
rect 425904 535394 426504 571158
rect 425904 535158 426086 535394
rect 426322 535158 426504 535394
rect 425904 499394 426504 535158
rect 425904 499158 426086 499394
rect 426322 499158 426504 499394
rect 425904 463394 426504 499158
rect 425904 463158 426086 463394
rect 426322 463158 426504 463394
rect 425904 427394 426504 463158
rect 425904 427158 426086 427394
rect 426322 427158 426504 427394
rect 425904 425308 426504 427158
rect 432804 704838 433404 705830
rect 432804 704602 432986 704838
rect 433222 704602 433404 704838
rect 432804 704518 433404 704602
rect 432804 704282 432986 704518
rect 433222 704282 433404 704518
rect 432804 686294 433404 704282
rect 432804 686058 432986 686294
rect 433222 686058 433404 686294
rect 432804 650294 433404 686058
rect 432804 650058 432986 650294
rect 433222 650058 433404 650294
rect 432804 614294 433404 650058
rect 432804 614058 432986 614294
rect 433222 614058 433404 614294
rect 432804 578294 433404 614058
rect 432804 578058 432986 578294
rect 433222 578058 433404 578294
rect 432804 542294 433404 578058
rect 432804 542058 432986 542294
rect 433222 542058 433404 542294
rect 432804 506294 433404 542058
rect 432804 506058 432986 506294
rect 433222 506058 433404 506294
rect 432804 470294 433404 506058
rect 432804 470058 432986 470294
rect 433222 470058 433404 470294
rect 432804 434294 433404 470058
rect 432804 434058 432986 434294
rect 433222 434058 433404 434294
rect 432804 425308 433404 434058
rect 436504 689994 437104 706202
rect 436504 689758 436686 689994
rect 436922 689758 437104 689994
rect 436504 653994 437104 689758
rect 436504 653758 436686 653994
rect 436922 653758 437104 653994
rect 436504 617994 437104 653758
rect 436504 617758 436686 617994
rect 436922 617758 437104 617994
rect 436504 581994 437104 617758
rect 436504 581758 436686 581994
rect 436922 581758 437104 581994
rect 436504 545994 437104 581758
rect 436504 545758 436686 545994
rect 436922 545758 437104 545994
rect 436504 509994 437104 545758
rect 436504 509758 436686 509994
rect 436922 509758 437104 509994
rect 436504 473994 437104 509758
rect 436504 473758 436686 473994
rect 436922 473758 437104 473994
rect 436504 437994 437104 473758
rect 436504 437758 436686 437994
rect 436922 437758 437104 437994
rect 436504 425308 437104 437758
rect 440204 693694 440804 708122
rect 440204 693458 440386 693694
rect 440622 693458 440804 693694
rect 440204 657694 440804 693458
rect 440204 657458 440386 657694
rect 440622 657458 440804 657694
rect 440204 621694 440804 657458
rect 440204 621458 440386 621694
rect 440622 621458 440804 621694
rect 440204 585694 440804 621458
rect 440204 585458 440386 585694
rect 440622 585458 440804 585694
rect 440204 549694 440804 585458
rect 440204 549458 440386 549694
rect 440622 549458 440804 549694
rect 440204 513694 440804 549458
rect 440204 513458 440386 513694
rect 440622 513458 440804 513694
rect 440204 477694 440804 513458
rect 440204 477458 440386 477694
rect 440622 477458 440804 477694
rect 440204 441694 440804 477458
rect 440204 441458 440386 441694
rect 440622 441458 440804 441694
rect 440204 425308 440804 441458
rect 443904 697394 444504 710042
rect 461904 711558 462504 711590
rect 461904 711322 462086 711558
rect 462322 711322 462504 711558
rect 461904 711238 462504 711322
rect 461904 711002 462086 711238
rect 462322 711002 462504 711238
rect 458204 709638 458804 709670
rect 458204 709402 458386 709638
rect 458622 709402 458804 709638
rect 458204 709318 458804 709402
rect 458204 709082 458386 709318
rect 458622 709082 458804 709318
rect 454504 707718 455104 707750
rect 454504 707482 454686 707718
rect 454922 707482 455104 707718
rect 454504 707398 455104 707482
rect 454504 707162 454686 707398
rect 454922 707162 455104 707398
rect 443904 697158 444086 697394
rect 444322 697158 444504 697394
rect 443904 661394 444504 697158
rect 443904 661158 444086 661394
rect 444322 661158 444504 661394
rect 443904 625394 444504 661158
rect 443904 625158 444086 625394
rect 444322 625158 444504 625394
rect 443904 589394 444504 625158
rect 443904 589158 444086 589394
rect 444322 589158 444504 589394
rect 443904 553394 444504 589158
rect 443904 553158 444086 553394
rect 444322 553158 444504 553394
rect 443904 517394 444504 553158
rect 443904 517158 444086 517394
rect 444322 517158 444504 517394
rect 443904 481394 444504 517158
rect 443904 481158 444086 481394
rect 444322 481158 444504 481394
rect 443904 445394 444504 481158
rect 443904 445158 444086 445394
rect 444322 445158 444504 445394
rect 443904 425308 444504 445158
rect 450804 705798 451404 705830
rect 450804 705562 450986 705798
rect 451222 705562 451404 705798
rect 450804 705478 451404 705562
rect 450804 705242 450986 705478
rect 451222 705242 451404 705478
rect 450804 668294 451404 705242
rect 450804 668058 450986 668294
rect 451222 668058 451404 668294
rect 450804 632294 451404 668058
rect 450804 632058 450986 632294
rect 451222 632058 451404 632294
rect 450804 596294 451404 632058
rect 450804 596058 450986 596294
rect 451222 596058 451404 596294
rect 450804 560294 451404 596058
rect 450804 560058 450986 560294
rect 451222 560058 451404 560294
rect 450804 524294 451404 560058
rect 450804 524058 450986 524294
rect 451222 524058 451404 524294
rect 450804 488294 451404 524058
rect 450804 488058 450986 488294
rect 451222 488058 451404 488294
rect 450804 452294 451404 488058
rect 450804 452058 450986 452294
rect 451222 452058 451404 452294
rect 450804 425308 451404 452058
rect 454504 671994 455104 707162
rect 454504 671758 454686 671994
rect 454922 671758 455104 671994
rect 454504 635994 455104 671758
rect 454504 635758 454686 635994
rect 454922 635758 455104 635994
rect 454504 599994 455104 635758
rect 454504 599758 454686 599994
rect 454922 599758 455104 599994
rect 454504 563994 455104 599758
rect 454504 563758 454686 563994
rect 454922 563758 455104 563994
rect 454504 527994 455104 563758
rect 454504 527758 454686 527994
rect 454922 527758 455104 527994
rect 454504 491994 455104 527758
rect 454504 491758 454686 491994
rect 454922 491758 455104 491994
rect 454504 455994 455104 491758
rect 454504 455758 454686 455994
rect 454922 455758 455104 455994
rect 454504 425308 455104 455758
rect 458204 675694 458804 709082
rect 458204 675458 458386 675694
rect 458622 675458 458804 675694
rect 458204 639694 458804 675458
rect 458204 639458 458386 639694
rect 458622 639458 458804 639694
rect 458204 603694 458804 639458
rect 458204 603458 458386 603694
rect 458622 603458 458804 603694
rect 458204 567694 458804 603458
rect 458204 567458 458386 567694
rect 458622 567458 458804 567694
rect 458204 531694 458804 567458
rect 458204 531458 458386 531694
rect 458622 531458 458804 531694
rect 458204 495694 458804 531458
rect 458204 495458 458386 495694
rect 458622 495458 458804 495694
rect 458204 459694 458804 495458
rect 458204 459458 458386 459694
rect 458622 459458 458804 459694
rect 458204 425308 458804 459458
rect 461904 679394 462504 711002
rect 479904 710598 480504 711590
rect 479904 710362 480086 710598
rect 480322 710362 480504 710598
rect 479904 710278 480504 710362
rect 479904 710042 480086 710278
rect 480322 710042 480504 710278
rect 476204 708678 476804 709670
rect 476204 708442 476386 708678
rect 476622 708442 476804 708678
rect 476204 708358 476804 708442
rect 476204 708122 476386 708358
rect 476622 708122 476804 708358
rect 472504 706758 473104 707750
rect 472504 706522 472686 706758
rect 472922 706522 473104 706758
rect 472504 706438 473104 706522
rect 472504 706202 472686 706438
rect 472922 706202 473104 706438
rect 461904 679158 462086 679394
rect 462322 679158 462504 679394
rect 461904 643394 462504 679158
rect 461904 643158 462086 643394
rect 462322 643158 462504 643394
rect 461904 607394 462504 643158
rect 461904 607158 462086 607394
rect 462322 607158 462504 607394
rect 461904 571394 462504 607158
rect 461904 571158 462086 571394
rect 462322 571158 462504 571394
rect 461904 535394 462504 571158
rect 461904 535158 462086 535394
rect 462322 535158 462504 535394
rect 461904 499394 462504 535158
rect 461904 499158 462086 499394
rect 462322 499158 462504 499394
rect 461904 463394 462504 499158
rect 461904 463158 462086 463394
rect 462322 463158 462504 463394
rect 461904 427394 462504 463158
rect 461904 427158 462086 427394
rect 462322 427158 462504 427394
rect 461904 425308 462504 427158
rect 468804 704838 469404 705830
rect 468804 704602 468986 704838
rect 469222 704602 469404 704838
rect 468804 704518 469404 704602
rect 468804 704282 468986 704518
rect 469222 704282 469404 704518
rect 468804 686294 469404 704282
rect 468804 686058 468986 686294
rect 469222 686058 469404 686294
rect 468804 650294 469404 686058
rect 468804 650058 468986 650294
rect 469222 650058 469404 650294
rect 468804 614294 469404 650058
rect 468804 614058 468986 614294
rect 469222 614058 469404 614294
rect 468804 578294 469404 614058
rect 468804 578058 468986 578294
rect 469222 578058 469404 578294
rect 468804 542294 469404 578058
rect 468804 542058 468986 542294
rect 469222 542058 469404 542294
rect 468804 506294 469404 542058
rect 468804 506058 468986 506294
rect 469222 506058 469404 506294
rect 468804 470294 469404 506058
rect 468804 470058 468986 470294
rect 469222 470058 469404 470294
rect 468804 434294 469404 470058
rect 468804 434058 468986 434294
rect 469222 434058 469404 434294
rect 468804 425308 469404 434058
rect 472504 689994 473104 706202
rect 472504 689758 472686 689994
rect 472922 689758 473104 689994
rect 472504 653994 473104 689758
rect 472504 653758 472686 653994
rect 472922 653758 473104 653994
rect 472504 617994 473104 653758
rect 472504 617758 472686 617994
rect 472922 617758 473104 617994
rect 472504 581994 473104 617758
rect 472504 581758 472686 581994
rect 472922 581758 473104 581994
rect 472504 545994 473104 581758
rect 472504 545758 472686 545994
rect 472922 545758 473104 545994
rect 472504 509994 473104 545758
rect 472504 509758 472686 509994
rect 472922 509758 473104 509994
rect 472504 473994 473104 509758
rect 472504 473758 472686 473994
rect 472922 473758 473104 473994
rect 472504 437994 473104 473758
rect 472504 437758 472686 437994
rect 472922 437758 473104 437994
rect 472504 425308 473104 437758
rect 476204 693694 476804 708122
rect 476204 693458 476386 693694
rect 476622 693458 476804 693694
rect 476204 657694 476804 693458
rect 476204 657458 476386 657694
rect 476622 657458 476804 657694
rect 476204 621694 476804 657458
rect 476204 621458 476386 621694
rect 476622 621458 476804 621694
rect 476204 585694 476804 621458
rect 476204 585458 476386 585694
rect 476622 585458 476804 585694
rect 476204 549694 476804 585458
rect 476204 549458 476386 549694
rect 476622 549458 476804 549694
rect 476204 513694 476804 549458
rect 476204 513458 476386 513694
rect 476622 513458 476804 513694
rect 476204 477694 476804 513458
rect 476204 477458 476386 477694
rect 476622 477458 476804 477694
rect 476204 441694 476804 477458
rect 476204 441458 476386 441694
rect 476622 441458 476804 441694
rect 476204 425308 476804 441458
rect 479904 697394 480504 710042
rect 497904 711558 498504 711590
rect 497904 711322 498086 711558
rect 498322 711322 498504 711558
rect 497904 711238 498504 711322
rect 497904 711002 498086 711238
rect 498322 711002 498504 711238
rect 494204 709638 494804 709670
rect 494204 709402 494386 709638
rect 494622 709402 494804 709638
rect 494204 709318 494804 709402
rect 494204 709082 494386 709318
rect 494622 709082 494804 709318
rect 490504 707718 491104 707750
rect 490504 707482 490686 707718
rect 490922 707482 491104 707718
rect 490504 707398 491104 707482
rect 490504 707162 490686 707398
rect 490922 707162 491104 707398
rect 479904 697158 480086 697394
rect 480322 697158 480504 697394
rect 479904 661394 480504 697158
rect 479904 661158 480086 661394
rect 480322 661158 480504 661394
rect 479904 625394 480504 661158
rect 479904 625158 480086 625394
rect 480322 625158 480504 625394
rect 479904 589394 480504 625158
rect 479904 589158 480086 589394
rect 480322 589158 480504 589394
rect 479904 553394 480504 589158
rect 479904 553158 480086 553394
rect 480322 553158 480504 553394
rect 479904 517394 480504 553158
rect 479904 517158 480086 517394
rect 480322 517158 480504 517394
rect 479904 481394 480504 517158
rect 479904 481158 480086 481394
rect 480322 481158 480504 481394
rect 479904 445394 480504 481158
rect 479904 445158 480086 445394
rect 480322 445158 480504 445394
rect 340272 416294 340620 416476
rect 340272 416058 340328 416294
rect 340564 416058 340620 416294
rect 340272 415876 340620 416058
rect 476000 416294 476348 416476
rect 476000 416058 476056 416294
rect 476292 416058 476348 416294
rect 476000 415876 476348 416058
rect 335904 409158 336086 409394
rect 336322 409158 336504 409394
rect 335904 373394 336504 409158
rect 479904 409394 480504 445158
rect 479904 409158 480086 409394
rect 480322 409158 480504 409394
rect 340952 398294 341300 398476
rect 340952 398058 341008 398294
rect 341244 398058 341300 398294
rect 340952 397876 341300 398058
rect 475320 398294 475668 398476
rect 475320 398058 475376 398294
rect 475612 398058 475668 398294
rect 475320 397876 475668 398058
rect 340272 380294 340620 380476
rect 340272 380058 340328 380294
rect 340564 380058 340620 380294
rect 340272 379876 340620 380058
rect 476000 380294 476348 380476
rect 476000 380058 476056 380294
rect 476292 380058 476348 380294
rect 476000 379876 476348 380058
rect 335904 373158 336086 373394
rect 336322 373158 336504 373394
rect 335904 337394 336504 373158
rect 479904 373394 480504 409158
rect 479904 373158 480086 373394
rect 480322 373158 480504 373394
rect 340952 362294 341300 362476
rect 340952 362058 341008 362294
rect 341244 362058 341300 362294
rect 340952 361876 341300 362058
rect 475320 362294 475668 362476
rect 475320 362058 475376 362294
rect 475612 362058 475668 362294
rect 475320 361876 475668 362058
rect 340272 344294 340620 344476
rect 340272 344058 340328 344294
rect 340564 344058 340620 344294
rect 340272 343876 340620 344058
rect 476000 344294 476348 344476
rect 476000 344058 476056 344294
rect 476292 344058 476348 344294
rect 476000 343876 476348 344058
rect 356056 339690 356116 340000
rect 357144 339690 357204 340000
rect 358232 339690 358292 340000
rect 356056 339630 356162 339690
rect 356102 338061 356162 339630
rect 357022 339630 357204 339690
rect 358126 339630 358292 339690
rect 359592 339690 359652 340000
rect 360544 339690 360604 340000
rect 359592 339630 359658 339690
rect 356099 338060 356165 338061
rect 335904 337158 336086 337394
rect 336322 337158 336504 337394
rect 335904 301394 336504 337158
rect 335904 301158 336086 301394
rect 336322 301158 336504 301394
rect 335904 265394 336504 301158
rect 335904 265158 336086 265394
rect 336322 265158 336504 265394
rect 335904 229394 336504 265158
rect 335904 229158 336086 229394
rect 336322 229158 336504 229394
rect 335904 193394 336504 229158
rect 335904 193158 336086 193394
rect 336322 193158 336504 193394
rect 335904 157394 336504 193158
rect 335904 157158 336086 157394
rect 336322 157158 336504 157394
rect 335904 121394 336504 157158
rect 335904 121158 336086 121394
rect 336322 121158 336504 121394
rect 335904 85394 336504 121158
rect 335904 85158 336086 85394
rect 336322 85158 336504 85394
rect 335904 49394 336504 85158
rect 335904 49158 336086 49394
rect 336322 49158 336504 49394
rect 335904 13394 336504 49158
rect 335904 13158 336086 13394
rect 336322 13158 336504 13394
rect 317904 -7302 318086 -7066
rect 318322 -7302 318504 -7066
rect 317904 -7386 318504 -7302
rect 317904 -7622 318086 -7386
rect 318322 -7622 318504 -7386
rect 317904 -7654 318504 -7622
rect 335904 -6106 336504 13158
rect 342804 308294 343404 338000
rect 342804 308058 342986 308294
rect 343222 308058 343404 308294
rect 342804 272294 343404 308058
rect 342804 272058 342986 272294
rect 343222 272058 343404 272294
rect 342804 236294 343404 272058
rect 342804 236058 342986 236294
rect 343222 236058 343404 236294
rect 342804 200294 343404 236058
rect 342804 200058 342986 200294
rect 343222 200058 343404 200294
rect 342804 164294 343404 200058
rect 342804 164058 342986 164294
rect 343222 164058 343404 164294
rect 342804 128294 343404 164058
rect 342804 128058 342986 128294
rect 343222 128058 343404 128294
rect 342804 92294 343404 128058
rect 342804 92058 342986 92294
rect 343222 92058 343404 92294
rect 342804 56294 343404 92058
rect 342804 56058 342986 56294
rect 343222 56058 343404 56294
rect 342804 20294 343404 56058
rect 342804 20058 342986 20294
rect 343222 20058 343404 20294
rect 342804 -1306 343404 20058
rect 342804 -1542 342986 -1306
rect 343222 -1542 343404 -1306
rect 342804 -1626 343404 -1542
rect 342804 -1862 342986 -1626
rect 343222 -1862 343404 -1626
rect 342804 -1894 343404 -1862
rect 346504 311994 347104 338000
rect 346504 311758 346686 311994
rect 346922 311758 347104 311994
rect 346504 275994 347104 311758
rect 346504 275758 346686 275994
rect 346922 275758 347104 275994
rect 346504 239994 347104 275758
rect 346504 239758 346686 239994
rect 346922 239758 347104 239994
rect 346504 203994 347104 239758
rect 346504 203758 346686 203994
rect 346922 203758 347104 203994
rect 346504 167994 347104 203758
rect 346504 167758 346686 167994
rect 346922 167758 347104 167994
rect 346504 131994 347104 167758
rect 346504 131758 346686 131994
rect 346922 131758 347104 131994
rect 346504 95994 347104 131758
rect 346504 95758 346686 95994
rect 346922 95758 347104 95994
rect 346504 59994 347104 95758
rect 346504 59758 346686 59994
rect 346922 59758 347104 59994
rect 346504 23994 347104 59758
rect 346504 23758 346686 23994
rect 346922 23758 347104 23994
rect 346504 -3226 347104 23758
rect 346504 -3462 346686 -3226
rect 346922 -3462 347104 -3226
rect 346504 -3546 347104 -3462
rect 346504 -3782 346686 -3546
rect 346922 -3782 347104 -3546
rect 346504 -3814 347104 -3782
rect 350204 315694 350804 338000
rect 350204 315458 350386 315694
rect 350622 315458 350804 315694
rect 350204 279694 350804 315458
rect 350204 279458 350386 279694
rect 350622 279458 350804 279694
rect 350204 243694 350804 279458
rect 350204 243458 350386 243694
rect 350622 243458 350804 243694
rect 350204 207694 350804 243458
rect 350204 207458 350386 207694
rect 350622 207458 350804 207694
rect 350204 171694 350804 207458
rect 350204 171458 350386 171694
rect 350622 171458 350804 171694
rect 350204 135694 350804 171458
rect 350204 135458 350386 135694
rect 350622 135458 350804 135694
rect 350204 99694 350804 135458
rect 350204 99458 350386 99694
rect 350622 99458 350804 99694
rect 350204 63694 350804 99458
rect 350204 63458 350386 63694
rect 350622 63458 350804 63694
rect 350204 27694 350804 63458
rect 350204 27458 350386 27694
rect 350622 27458 350804 27694
rect 350204 -5146 350804 27458
rect 350204 -5382 350386 -5146
rect 350622 -5382 350804 -5146
rect 350204 -5466 350804 -5382
rect 350204 -5702 350386 -5466
rect 350622 -5702 350804 -5466
rect 350204 -5734 350804 -5702
rect 353904 319394 354504 338000
rect 356099 337996 356100 338060
rect 356164 337996 356165 338060
rect 356099 337995 356165 337996
rect 357022 337653 357082 339630
rect 358126 337653 358186 339630
rect 359598 337653 359658 339630
rect 360518 339630 360604 339690
rect 361768 339690 361828 340000
rect 363128 339690 363188 340000
rect 364216 339690 364276 340000
rect 361768 339630 361866 339690
rect 360518 337653 360578 339630
rect 357019 337652 357085 337653
rect 357019 337588 357020 337652
rect 357084 337588 357085 337652
rect 357019 337587 357085 337588
rect 358123 337652 358189 337653
rect 358123 337588 358124 337652
rect 358188 337588 358189 337652
rect 358123 337587 358189 337588
rect 359595 337652 359661 337653
rect 359595 337588 359596 337652
rect 359660 337588 359661 337652
rect 359595 337587 359661 337588
rect 360515 337652 360581 337653
rect 360515 337588 360516 337652
rect 360580 337588 360581 337652
rect 360515 337587 360581 337588
rect 353904 319158 354086 319394
rect 354322 319158 354504 319394
rect 353904 283394 354504 319158
rect 353904 283158 354086 283394
rect 354322 283158 354504 283394
rect 353904 247394 354504 283158
rect 353904 247158 354086 247394
rect 354322 247158 354504 247394
rect 353904 211394 354504 247158
rect 353904 211158 354086 211394
rect 354322 211158 354504 211394
rect 353904 175394 354504 211158
rect 353904 175158 354086 175394
rect 354322 175158 354504 175394
rect 353904 139394 354504 175158
rect 353904 139158 354086 139394
rect 354322 139158 354504 139394
rect 353904 103394 354504 139158
rect 353904 103158 354086 103394
rect 354322 103158 354504 103394
rect 353904 67394 354504 103158
rect 353904 67158 354086 67394
rect 354322 67158 354504 67394
rect 353904 31394 354504 67158
rect 353904 31158 354086 31394
rect 354322 31158 354504 31394
rect 335904 -6342 336086 -6106
rect 336322 -6342 336504 -6106
rect 335904 -6426 336504 -6342
rect 335904 -6662 336086 -6426
rect 336322 -6662 336504 -6426
rect 335904 -7654 336504 -6662
rect 353904 -7066 354504 31158
rect 360804 326294 361404 338000
rect 361806 337109 361866 339630
rect 363094 339630 363188 339690
rect 364198 339630 364276 339690
rect 363094 337653 363154 339630
rect 364198 337789 364258 339630
rect 365440 339510 365500 340000
rect 366528 339510 366588 340000
rect 367616 339510 367676 340000
rect 368296 339510 368356 340000
rect 365440 339450 365546 339510
rect 364195 337788 364261 337789
rect 364195 337724 364196 337788
rect 364260 337724 364261 337788
rect 364195 337723 364261 337724
rect 363091 337652 363157 337653
rect 363091 337588 363092 337652
rect 363156 337588 363157 337652
rect 363091 337587 363157 337588
rect 361803 337108 361869 337109
rect 361803 337044 361804 337108
rect 361868 337044 361869 337108
rect 361803 337043 361869 337044
rect 360804 326058 360986 326294
rect 361222 326058 361404 326294
rect 360804 290294 361404 326058
rect 360804 290058 360986 290294
rect 361222 290058 361404 290294
rect 360804 254294 361404 290058
rect 360804 254058 360986 254294
rect 361222 254058 361404 254294
rect 360804 218294 361404 254058
rect 360804 218058 360986 218294
rect 361222 218058 361404 218294
rect 360804 182294 361404 218058
rect 360804 182058 360986 182294
rect 361222 182058 361404 182294
rect 360804 146294 361404 182058
rect 360804 146058 360986 146294
rect 361222 146058 361404 146294
rect 360804 110294 361404 146058
rect 360804 110058 360986 110294
rect 361222 110058 361404 110294
rect 360804 74294 361404 110058
rect 360804 74058 360986 74294
rect 361222 74058 361404 74294
rect 360804 38294 361404 74058
rect 360804 38058 360986 38294
rect 361222 38058 361404 38294
rect 360804 2294 361404 38058
rect 360804 2058 360986 2294
rect 361222 2058 361404 2294
rect 360804 -346 361404 2058
rect 360804 -582 360986 -346
rect 361222 -582 361404 -346
rect 360804 -666 361404 -582
rect 360804 -902 360986 -666
rect 361222 -902 361404 -666
rect 360804 -1894 361404 -902
rect 364504 329994 365104 338000
rect 365486 337653 365546 339450
rect 366406 339450 366588 339510
rect 367510 339450 367676 339510
rect 368062 339450 368356 339510
rect 368704 339510 368764 340000
rect 370064 339510 370124 340000
rect 370744 339510 370804 340000
rect 368704 339450 369042 339510
rect 370064 339450 370146 339510
rect 366406 337653 366466 339450
rect 367510 337653 367570 339450
rect 368062 337789 368122 339450
rect 368982 338061 369042 339450
rect 368979 338060 369045 338061
rect 368059 337788 368125 337789
rect 368059 337724 368060 337788
rect 368124 337724 368125 337788
rect 368059 337723 368125 337724
rect 365483 337652 365549 337653
rect 365483 337588 365484 337652
rect 365548 337588 365549 337652
rect 365483 337587 365549 337588
rect 366403 337652 366469 337653
rect 366403 337588 366404 337652
rect 366468 337588 366469 337652
rect 366403 337587 366469 337588
rect 367507 337652 367573 337653
rect 367507 337588 367508 337652
rect 367572 337588 367573 337652
rect 367507 337587 367573 337588
rect 364504 329758 364686 329994
rect 364922 329758 365104 329994
rect 364504 293994 365104 329758
rect 364504 293758 364686 293994
rect 364922 293758 365104 293994
rect 364504 257994 365104 293758
rect 364504 257758 364686 257994
rect 364922 257758 365104 257994
rect 364504 221994 365104 257758
rect 364504 221758 364686 221994
rect 364922 221758 365104 221994
rect 364504 185994 365104 221758
rect 364504 185758 364686 185994
rect 364922 185758 365104 185994
rect 364504 149994 365104 185758
rect 364504 149758 364686 149994
rect 364922 149758 365104 149994
rect 364504 113994 365104 149758
rect 364504 113758 364686 113994
rect 364922 113758 365104 113994
rect 364504 77994 365104 113758
rect 364504 77758 364686 77994
rect 364922 77758 365104 77994
rect 364504 41994 365104 77758
rect 364504 41758 364686 41994
rect 364922 41758 365104 41994
rect 364504 5994 365104 41758
rect 364504 5758 364686 5994
rect 364922 5758 365104 5994
rect 364504 -2266 365104 5758
rect 364504 -2502 364686 -2266
rect 364922 -2502 365104 -2266
rect 364504 -2586 365104 -2502
rect 364504 -2822 364686 -2586
rect 364922 -2822 365104 -2586
rect 364504 -3814 365104 -2822
rect 368204 333694 368804 338000
rect 368979 337996 368980 338060
rect 369044 337996 369045 338060
rect 368979 337995 369045 337996
rect 370086 336973 370146 339450
rect 370638 339450 370804 339510
rect 371288 339510 371348 340000
rect 372376 339510 372436 340000
rect 373464 339690 373524 340000
rect 371288 339450 371434 339510
rect 370083 336972 370149 336973
rect 370083 336908 370084 336972
rect 370148 336908 370149 336972
rect 370083 336907 370149 336908
rect 370638 336837 370698 339450
rect 371374 337653 371434 339450
rect 372294 339450 372436 339510
rect 373398 339630 373524 339690
rect 372294 338197 372354 339450
rect 372291 338196 372357 338197
rect 372291 338132 372292 338196
rect 372356 338132 372357 338196
rect 372291 338131 372357 338132
rect 371371 337652 371437 337653
rect 371371 337588 371372 337652
rect 371436 337588 371437 337652
rect 371371 337587 371437 337588
rect 371904 337394 372504 338000
rect 373398 337653 373458 339630
rect 373600 339510 373660 340000
rect 374552 339510 374612 340000
rect 375912 339690 375972 340000
rect 373582 339450 373660 339510
rect 374502 339450 374612 339510
rect 375790 339630 375972 339690
rect 373582 337789 373642 339450
rect 373579 337788 373645 337789
rect 373579 337724 373580 337788
rect 373644 337724 373645 337788
rect 373579 337723 373645 337724
rect 374502 337653 374562 339450
rect 373395 337652 373461 337653
rect 373395 337588 373396 337652
rect 373460 337588 373461 337652
rect 373395 337587 373461 337588
rect 374499 337652 374565 337653
rect 374499 337588 374500 337652
rect 374564 337588 374565 337652
rect 374499 337587 374565 337588
rect 371904 337158 372086 337394
rect 372322 337158 372504 337394
rect 375790 337245 375850 339630
rect 376048 339510 376108 340000
rect 377000 339510 377060 340000
rect 378088 339510 378148 340000
rect 375974 339450 376108 339510
rect 376894 339450 377060 339510
rect 377998 339450 378148 339510
rect 378496 339510 378556 340000
rect 379448 339690 379508 340000
rect 379448 339630 379530 339690
rect 378496 339450 378610 339510
rect 375787 337244 375853 337245
rect 375787 337180 375788 337244
rect 375852 337180 375853 337244
rect 375787 337179 375853 337180
rect 370635 336836 370701 336837
rect 370635 336772 370636 336836
rect 370700 336772 370701 336836
rect 370635 336771 370701 336772
rect 368204 333458 368386 333694
rect 368622 333458 368804 333694
rect 368204 297694 368804 333458
rect 368204 297458 368386 297694
rect 368622 297458 368804 297694
rect 368204 261694 368804 297458
rect 368204 261458 368386 261694
rect 368622 261458 368804 261694
rect 368204 225694 368804 261458
rect 368204 225458 368386 225694
rect 368622 225458 368804 225694
rect 368204 189694 368804 225458
rect 368204 189458 368386 189694
rect 368622 189458 368804 189694
rect 368204 153694 368804 189458
rect 368204 153458 368386 153694
rect 368622 153458 368804 153694
rect 368204 117694 368804 153458
rect 368204 117458 368386 117694
rect 368622 117458 368804 117694
rect 368204 81694 368804 117458
rect 368204 81458 368386 81694
rect 368622 81458 368804 81694
rect 368204 45694 368804 81458
rect 368204 45458 368386 45694
rect 368622 45458 368804 45694
rect 368204 9694 368804 45458
rect 368204 9458 368386 9694
rect 368622 9458 368804 9694
rect 368204 -4186 368804 9458
rect 368204 -4422 368386 -4186
rect 368622 -4422 368804 -4186
rect 368204 -4506 368804 -4422
rect 368204 -4742 368386 -4506
rect 368622 -4742 368804 -4506
rect 368204 -5734 368804 -4742
rect 371904 301394 372504 337158
rect 375974 337109 376034 339450
rect 376894 337653 376954 339450
rect 377998 337789 378058 339450
rect 378550 337925 378610 339450
rect 378547 337924 378613 337925
rect 378547 337860 378548 337924
rect 378612 337860 378613 337924
rect 378547 337859 378613 337860
rect 377995 337788 378061 337789
rect 377995 337724 377996 337788
rect 378060 337724 378061 337788
rect 377995 337723 378061 337724
rect 376891 337652 376957 337653
rect 376891 337588 376892 337652
rect 376956 337588 376957 337652
rect 376891 337587 376957 337588
rect 375971 337108 376037 337109
rect 375971 337044 375972 337108
rect 376036 337044 376037 337108
rect 375971 337043 376037 337044
rect 371904 301158 372086 301394
rect 372322 301158 372504 301394
rect 371904 265394 372504 301158
rect 371904 265158 372086 265394
rect 372322 265158 372504 265394
rect 371904 229394 372504 265158
rect 371904 229158 372086 229394
rect 372322 229158 372504 229394
rect 371904 193394 372504 229158
rect 371904 193158 372086 193394
rect 372322 193158 372504 193394
rect 371904 157394 372504 193158
rect 371904 157158 372086 157394
rect 372322 157158 372504 157394
rect 371904 121394 372504 157158
rect 371904 121158 372086 121394
rect 372322 121158 372504 121394
rect 371904 85394 372504 121158
rect 371904 85158 372086 85394
rect 372322 85158 372504 85394
rect 371904 49394 372504 85158
rect 371904 49158 372086 49394
rect 372322 49158 372504 49394
rect 371904 13394 372504 49158
rect 371904 13158 372086 13394
rect 372322 13158 372504 13394
rect 353904 -7302 354086 -7066
rect 354322 -7302 354504 -7066
rect 353904 -7386 354504 -7302
rect 353904 -7622 354086 -7386
rect 354322 -7622 354504 -7386
rect 353904 -7654 354504 -7622
rect 371904 -6106 372504 13158
rect 378804 308294 379404 338000
rect 379470 337653 379530 339630
rect 380672 339510 380732 340000
rect 380574 339450 380732 339510
rect 381080 339510 381140 340000
rect 381760 339510 381820 340000
rect 382848 339510 382908 340000
rect 383528 339510 383588 340000
rect 383936 339510 383996 340000
rect 385296 339510 385356 340000
rect 385976 339510 386036 340000
rect 381080 339450 381186 339510
rect 380574 337789 380634 339450
rect 380571 337788 380637 337789
rect 380571 337724 380572 337788
rect 380636 337724 380637 337788
rect 380571 337723 380637 337724
rect 381126 337653 381186 339450
rect 381678 339450 381820 339510
rect 382782 339450 382908 339510
rect 383518 339450 383588 339510
rect 383886 339450 383996 339510
rect 385174 339450 385356 339510
rect 385910 339450 386036 339510
rect 386384 339510 386444 340000
rect 387608 339510 387668 340000
rect 386384 339450 386522 339510
rect 379467 337652 379533 337653
rect 379467 337588 379468 337652
rect 379532 337588 379533 337652
rect 379467 337587 379533 337588
rect 381123 337652 381189 337653
rect 381123 337588 381124 337652
rect 381188 337588 381189 337652
rect 381123 337587 381189 337588
rect 381678 337381 381738 339450
rect 382782 338197 382842 339450
rect 382779 338196 382845 338197
rect 382779 338132 382780 338196
rect 382844 338132 382845 338196
rect 382779 338131 382845 338132
rect 381675 337380 381741 337381
rect 381675 337316 381676 337380
rect 381740 337316 381741 337380
rect 381675 337315 381741 337316
rect 378804 308058 378986 308294
rect 379222 308058 379404 308294
rect 378804 272294 379404 308058
rect 378804 272058 378986 272294
rect 379222 272058 379404 272294
rect 378804 236294 379404 272058
rect 378804 236058 378986 236294
rect 379222 236058 379404 236294
rect 378804 200294 379404 236058
rect 378804 200058 378986 200294
rect 379222 200058 379404 200294
rect 378804 164294 379404 200058
rect 378804 164058 378986 164294
rect 379222 164058 379404 164294
rect 378804 128294 379404 164058
rect 378804 128058 378986 128294
rect 379222 128058 379404 128294
rect 378804 92294 379404 128058
rect 378804 92058 378986 92294
rect 379222 92058 379404 92294
rect 378804 56294 379404 92058
rect 378804 56058 378986 56294
rect 379222 56058 379404 56294
rect 378804 20294 379404 56058
rect 378804 20058 378986 20294
rect 379222 20058 379404 20294
rect 378804 -1306 379404 20058
rect 378804 -1542 378986 -1306
rect 379222 -1542 379404 -1306
rect 378804 -1626 379404 -1542
rect 378804 -1862 378986 -1626
rect 379222 -1862 379404 -1626
rect 378804 -1894 379404 -1862
rect 382504 311994 383104 338000
rect 383518 337245 383578 339450
rect 383886 337653 383946 339450
rect 385174 337653 385234 339450
rect 383883 337652 383949 337653
rect 383883 337588 383884 337652
rect 383948 337588 383949 337652
rect 383883 337587 383949 337588
rect 385171 337652 385237 337653
rect 385171 337588 385172 337652
rect 385236 337588 385237 337652
rect 385171 337587 385237 337588
rect 383515 337244 383581 337245
rect 383515 337180 383516 337244
rect 383580 337180 383581 337244
rect 383515 337179 383581 337180
rect 385910 337109 385970 339450
rect 386462 338197 386522 339450
rect 387566 339450 387668 339510
rect 388288 339510 388348 340000
rect 388696 339510 388756 340000
rect 389784 339510 389844 340000
rect 391008 339690 391068 340000
rect 388288 339450 388362 339510
rect 386459 338196 386525 338197
rect 386459 338132 386460 338196
rect 386524 338132 386525 338196
rect 386459 338131 386525 338132
rect 385907 337108 385973 337109
rect 385907 337044 385908 337108
rect 385972 337044 385973 337108
rect 385907 337043 385973 337044
rect 382504 311758 382686 311994
rect 382922 311758 383104 311994
rect 382504 275994 383104 311758
rect 382504 275758 382686 275994
rect 382922 275758 383104 275994
rect 382504 239994 383104 275758
rect 382504 239758 382686 239994
rect 382922 239758 383104 239994
rect 382504 203994 383104 239758
rect 382504 203758 382686 203994
rect 382922 203758 383104 203994
rect 382504 167994 383104 203758
rect 382504 167758 382686 167994
rect 382922 167758 383104 167994
rect 382504 131994 383104 167758
rect 382504 131758 382686 131994
rect 382922 131758 383104 131994
rect 382504 95994 383104 131758
rect 382504 95758 382686 95994
rect 382922 95758 383104 95994
rect 382504 59994 383104 95758
rect 382504 59758 382686 59994
rect 382922 59758 383104 59994
rect 382504 23994 383104 59758
rect 382504 23758 382686 23994
rect 382922 23758 383104 23994
rect 382504 -3226 383104 23758
rect 382504 -3462 382686 -3226
rect 382922 -3462 383104 -3226
rect 382504 -3546 383104 -3462
rect 382504 -3782 382686 -3546
rect 382922 -3782 383104 -3546
rect 382504 -3814 383104 -3782
rect 386204 315694 386804 338000
rect 387566 337653 387626 339450
rect 388302 337653 388362 339450
rect 388670 339450 388756 339510
rect 389774 339450 389844 339510
rect 390878 339630 391068 339690
rect 388670 337789 388730 339450
rect 388667 337788 388733 337789
rect 388667 337724 388668 337788
rect 388732 337724 388733 337788
rect 388667 337723 388733 337724
rect 389774 337653 389834 339450
rect 387563 337652 387629 337653
rect 387563 337588 387564 337652
rect 387628 337588 387629 337652
rect 387563 337587 387629 337588
rect 388299 337652 388365 337653
rect 388299 337588 388300 337652
rect 388364 337588 388365 337652
rect 388299 337587 388365 337588
rect 389771 337652 389837 337653
rect 389771 337588 389772 337652
rect 389836 337588 389837 337652
rect 389771 337587 389837 337588
rect 386204 315458 386386 315694
rect 386622 315458 386804 315694
rect 386204 279694 386804 315458
rect 386204 279458 386386 279694
rect 386622 279458 386804 279694
rect 386204 243694 386804 279458
rect 386204 243458 386386 243694
rect 386622 243458 386804 243694
rect 386204 207694 386804 243458
rect 386204 207458 386386 207694
rect 386622 207458 386804 207694
rect 386204 171694 386804 207458
rect 386204 171458 386386 171694
rect 386622 171458 386804 171694
rect 386204 135694 386804 171458
rect 386204 135458 386386 135694
rect 386622 135458 386804 135694
rect 386204 99694 386804 135458
rect 386204 99458 386386 99694
rect 386622 99458 386804 99694
rect 386204 63694 386804 99458
rect 386204 63458 386386 63694
rect 386622 63458 386804 63694
rect 386204 27694 386804 63458
rect 386204 27458 386386 27694
rect 386622 27458 386804 27694
rect 386204 -5146 386804 27458
rect 386204 -5382 386386 -5146
rect 386622 -5382 386804 -5146
rect 386204 -5466 386804 -5382
rect 386204 -5702 386386 -5466
rect 386622 -5702 386804 -5466
rect 386204 -5734 386804 -5702
rect 389904 319394 390504 338000
rect 390878 337517 390938 339630
rect 391144 339510 391204 340000
rect 392232 339510 392292 340000
rect 391062 339450 391204 339510
rect 392166 339450 392292 339510
rect 391062 337789 391122 339450
rect 392166 337925 392226 339450
rect 393320 339010 393380 340000
rect 393592 339690 393652 340000
rect 394408 339690 394468 340000
rect 395768 339690 395828 340000
rect 396040 339690 396100 340000
rect 396992 339690 397052 340000
rect 398080 339690 398140 340000
rect 398488 339690 398548 340000
rect 399168 339690 399228 340000
rect 393592 339630 393698 339690
rect 393320 338950 393514 339010
rect 392163 337924 392229 337925
rect 392163 337860 392164 337924
rect 392228 337860 392229 337924
rect 392163 337859 392229 337860
rect 391059 337788 391125 337789
rect 391059 337724 391060 337788
rect 391124 337724 391125 337788
rect 391059 337723 391125 337724
rect 390875 337516 390941 337517
rect 390875 337452 390876 337516
rect 390940 337452 390941 337516
rect 390875 337451 390941 337452
rect 393454 336973 393514 338950
rect 393638 337653 393698 339630
rect 394374 339630 394468 339690
rect 395662 339630 395828 339690
rect 396030 339630 396100 339690
rect 396582 339630 397052 339690
rect 398054 339630 398140 339690
rect 398422 339630 398548 339690
rect 399158 339630 399228 339690
rect 400936 339690 400996 340000
rect 403520 339690 403580 340000
rect 405968 339690 406028 340000
rect 408280 339690 408340 340000
rect 411000 339690 411060 340000
rect 413448 339690 413508 340000
rect 400936 339630 401242 339690
rect 403520 339630 403634 339690
rect 393635 337652 393701 337653
rect 393635 337588 393636 337652
rect 393700 337588 393701 337652
rect 393635 337587 393701 337588
rect 394374 337517 394434 339630
rect 395662 337925 395722 339630
rect 395659 337924 395725 337925
rect 395659 337860 395660 337924
rect 395724 337860 395725 337924
rect 395659 337859 395725 337860
rect 396030 337653 396090 339630
rect 396582 337925 396642 339630
rect 396579 337924 396645 337925
rect 396579 337860 396580 337924
rect 396644 337860 396645 337924
rect 396579 337859 396645 337860
rect 396027 337652 396093 337653
rect 396027 337588 396028 337652
rect 396092 337588 396093 337652
rect 396027 337587 396093 337588
rect 394371 337516 394437 337517
rect 394371 337452 394372 337516
rect 394436 337452 394437 337516
rect 394371 337451 394437 337452
rect 393451 336972 393517 336973
rect 393451 336908 393452 336972
rect 393516 336908 393517 336972
rect 393451 336907 393517 336908
rect 389904 319158 390086 319394
rect 390322 319158 390504 319394
rect 389904 283394 390504 319158
rect 389904 283158 390086 283394
rect 390322 283158 390504 283394
rect 389904 247394 390504 283158
rect 389904 247158 390086 247394
rect 390322 247158 390504 247394
rect 389904 211394 390504 247158
rect 389904 211158 390086 211394
rect 390322 211158 390504 211394
rect 389904 175394 390504 211158
rect 389904 175158 390086 175394
rect 390322 175158 390504 175394
rect 389904 139394 390504 175158
rect 389904 139158 390086 139394
rect 390322 139158 390504 139394
rect 389904 103394 390504 139158
rect 389904 103158 390086 103394
rect 390322 103158 390504 103394
rect 389904 67394 390504 103158
rect 389904 67158 390086 67394
rect 390322 67158 390504 67394
rect 389904 31394 390504 67158
rect 389904 31158 390086 31394
rect 390322 31158 390504 31394
rect 371904 -6342 372086 -6106
rect 372322 -6342 372504 -6106
rect 371904 -6426 372504 -6342
rect 371904 -6662 372086 -6426
rect 372322 -6662 372504 -6426
rect 371904 -7654 372504 -6662
rect 389904 -7066 390504 31158
rect 396804 326294 397404 338000
rect 398054 337381 398114 339630
rect 398422 337653 398482 339630
rect 399158 337925 399218 339630
rect 399155 337924 399221 337925
rect 399155 337860 399156 337924
rect 399220 337860 399221 337924
rect 399155 337859 399221 337860
rect 398419 337652 398485 337653
rect 398419 337588 398420 337652
rect 398484 337588 398485 337652
rect 398419 337587 398485 337588
rect 398051 337380 398117 337381
rect 398051 337316 398052 337380
rect 398116 337316 398117 337380
rect 398051 337315 398117 337316
rect 396804 326058 396986 326294
rect 397222 326058 397404 326294
rect 396804 290294 397404 326058
rect 396804 290058 396986 290294
rect 397222 290058 397404 290294
rect 396804 254294 397404 290058
rect 396804 254058 396986 254294
rect 397222 254058 397404 254294
rect 396804 218294 397404 254058
rect 396804 218058 396986 218294
rect 397222 218058 397404 218294
rect 396804 182294 397404 218058
rect 396804 182058 396986 182294
rect 397222 182058 397404 182294
rect 396804 146294 397404 182058
rect 396804 146058 396986 146294
rect 397222 146058 397404 146294
rect 396804 110294 397404 146058
rect 396804 110058 396986 110294
rect 397222 110058 397404 110294
rect 396804 74294 397404 110058
rect 396804 74058 396986 74294
rect 397222 74058 397404 74294
rect 396804 38294 397404 74058
rect 396804 38058 396986 38294
rect 397222 38058 397404 38294
rect 396804 2294 397404 38058
rect 396804 2058 396986 2294
rect 397222 2058 397404 2294
rect 396804 -346 397404 2058
rect 396804 -582 396986 -346
rect 397222 -582 397404 -346
rect 396804 -666 397404 -582
rect 396804 -902 396986 -666
rect 397222 -902 397404 -666
rect 396804 -1894 397404 -902
rect 400504 329994 401104 338000
rect 401182 336837 401242 339630
rect 403574 337653 403634 339630
rect 405966 339630 406028 339690
rect 408174 339630 408340 339690
rect 410934 339630 411060 339690
rect 413326 339630 413508 339690
rect 415896 339690 415956 340000
rect 418480 339690 418540 340000
rect 420928 339690 420988 340000
rect 423512 339690 423572 340000
rect 425960 339690 426020 340000
rect 415896 339630 415962 339690
rect 403571 337652 403637 337653
rect 403571 337588 403572 337652
rect 403636 337588 403637 337652
rect 403571 337587 403637 337588
rect 401179 336836 401245 336837
rect 401179 336772 401180 336836
rect 401244 336772 401245 336836
rect 401179 336771 401245 336772
rect 400504 329758 400686 329994
rect 400922 329758 401104 329994
rect 400504 293994 401104 329758
rect 400504 293758 400686 293994
rect 400922 293758 401104 293994
rect 400504 257994 401104 293758
rect 400504 257758 400686 257994
rect 400922 257758 401104 257994
rect 400504 221994 401104 257758
rect 400504 221758 400686 221994
rect 400922 221758 401104 221994
rect 400504 185994 401104 221758
rect 400504 185758 400686 185994
rect 400922 185758 401104 185994
rect 400504 149994 401104 185758
rect 400504 149758 400686 149994
rect 400922 149758 401104 149994
rect 400504 113994 401104 149758
rect 400504 113758 400686 113994
rect 400922 113758 401104 113994
rect 400504 77994 401104 113758
rect 400504 77758 400686 77994
rect 400922 77758 401104 77994
rect 400504 41994 401104 77758
rect 400504 41758 400686 41994
rect 400922 41758 401104 41994
rect 400504 5994 401104 41758
rect 400504 5758 400686 5994
rect 400922 5758 401104 5994
rect 400504 -2266 401104 5758
rect 400504 -2502 400686 -2266
rect 400922 -2502 401104 -2266
rect 400504 -2586 401104 -2502
rect 400504 -2822 400686 -2586
rect 400922 -2822 401104 -2586
rect 400504 -3814 401104 -2822
rect 404204 333694 404804 338000
rect 405966 337653 406026 339630
rect 408174 338197 408234 339630
rect 408171 338196 408237 338197
rect 408171 338132 408172 338196
rect 408236 338132 408237 338196
rect 408171 338131 408237 338132
rect 405963 337652 406029 337653
rect 405963 337588 405964 337652
rect 406028 337588 406029 337652
rect 405963 337587 406029 337588
rect 404204 333458 404386 333694
rect 404622 333458 404804 333694
rect 404204 297694 404804 333458
rect 404204 297458 404386 297694
rect 404622 297458 404804 297694
rect 404204 261694 404804 297458
rect 404204 261458 404386 261694
rect 404622 261458 404804 261694
rect 404204 225694 404804 261458
rect 404204 225458 404386 225694
rect 404622 225458 404804 225694
rect 404204 189694 404804 225458
rect 404204 189458 404386 189694
rect 404622 189458 404804 189694
rect 404204 153694 404804 189458
rect 404204 153458 404386 153694
rect 404622 153458 404804 153694
rect 404204 117694 404804 153458
rect 404204 117458 404386 117694
rect 404622 117458 404804 117694
rect 404204 81694 404804 117458
rect 404204 81458 404386 81694
rect 404622 81458 404804 81694
rect 404204 45694 404804 81458
rect 404204 45458 404386 45694
rect 404622 45458 404804 45694
rect 404204 9694 404804 45458
rect 404204 9458 404386 9694
rect 404622 9458 404804 9694
rect 404204 -4186 404804 9458
rect 404204 -4422 404386 -4186
rect 404622 -4422 404804 -4186
rect 404204 -4506 404804 -4422
rect 404204 -4742 404386 -4506
rect 404622 -4742 404804 -4506
rect 404204 -5734 404804 -4742
rect 407904 337394 408504 338000
rect 410934 337653 410994 339630
rect 413326 337653 413386 339630
rect 410931 337652 410997 337653
rect 410931 337588 410932 337652
rect 410996 337588 410997 337652
rect 410931 337587 410997 337588
rect 413323 337652 413389 337653
rect 413323 337588 413324 337652
rect 413388 337588 413389 337652
rect 413323 337587 413389 337588
rect 407904 337158 408086 337394
rect 408322 337158 408504 337394
rect 407904 301394 408504 337158
rect 407904 301158 408086 301394
rect 408322 301158 408504 301394
rect 407904 265394 408504 301158
rect 407904 265158 408086 265394
rect 408322 265158 408504 265394
rect 407904 229394 408504 265158
rect 407904 229158 408086 229394
rect 408322 229158 408504 229394
rect 407904 193394 408504 229158
rect 407904 193158 408086 193394
rect 408322 193158 408504 193394
rect 407904 157394 408504 193158
rect 407904 157158 408086 157394
rect 408322 157158 408504 157394
rect 407904 121394 408504 157158
rect 407904 121158 408086 121394
rect 408322 121158 408504 121394
rect 407904 85394 408504 121158
rect 407904 85158 408086 85394
rect 408322 85158 408504 85394
rect 407904 49394 408504 85158
rect 407904 49158 408086 49394
rect 408322 49158 408504 49394
rect 407904 13394 408504 49158
rect 407904 13158 408086 13394
rect 408322 13158 408504 13394
rect 389904 -7302 390086 -7066
rect 390322 -7302 390504 -7066
rect 389904 -7386 390504 -7302
rect 389904 -7622 390086 -7386
rect 390322 -7622 390504 -7386
rect 389904 -7654 390504 -7622
rect 407904 -6106 408504 13158
rect 414804 308294 415404 338000
rect 415902 337653 415962 339630
rect 418294 339630 418540 339690
rect 420870 339630 420988 339690
rect 423446 339630 423572 339690
rect 425654 339630 426020 339690
rect 428544 339690 428604 340000
rect 430992 339690 431052 340000
rect 428544 339630 428658 339690
rect 418294 337653 418354 339630
rect 415899 337652 415965 337653
rect 415899 337588 415900 337652
rect 415964 337588 415965 337652
rect 415899 337587 415965 337588
rect 418291 337652 418357 337653
rect 418291 337588 418292 337652
rect 418356 337588 418357 337652
rect 418291 337587 418357 337588
rect 414804 308058 414986 308294
rect 415222 308058 415404 308294
rect 414804 272294 415404 308058
rect 414804 272058 414986 272294
rect 415222 272058 415404 272294
rect 414804 236294 415404 272058
rect 414804 236058 414986 236294
rect 415222 236058 415404 236294
rect 414804 200294 415404 236058
rect 414804 200058 414986 200294
rect 415222 200058 415404 200294
rect 414804 164294 415404 200058
rect 414804 164058 414986 164294
rect 415222 164058 415404 164294
rect 414804 128294 415404 164058
rect 414804 128058 414986 128294
rect 415222 128058 415404 128294
rect 414804 92294 415404 128058
rect 414804 92058 414986 92294
rect 415222 92058 415404 92294
rect 414804 56294 415404 92058
rect 414804 56058 414986 56294
rect 415222 56058 415404 56294
rect 414804 20294 415404 56058
rect 414804 20058 414986 20294
rect 415222 20058 415404 20294
rect 414804 -1306 415404 20058
rect 414804 -1542 414986 -1306
rect 415222 -1542 415404 -1306
rect 414804 -1626 415404 -1542
rect 414804 -1862 414986 -1626
rect 415222 -1862 415404 -1626
rect 414804 -1894 415404 -1862
rect 418504 311994 419104 338000
rect 420870 337653 420930 339630
rect 420867 337652 420933 337653
rect 420867 337588 420868 337652
rect 420932 337588 420933 337652
rect 420867 337587 420933 337588
rect 418504 311758 418686 311994
rect 418922 311758 419104 311994
rect 418504 275994 419104 311758
rect 418504 275758 418686 275994
rect 418922 275758 419104 275994
rect 418504 239994 419104 275758
rect 418504 239758 418686 239994
rect 418922 239758 419104 239994
rect 418504 203994 419104 239758
rect 418504 203758 418686 203994
rect 418922 203758 419104 203994
rect 418504 167994 419104 203758
rect 418504 167758 418686 167994
rect 418922 167758 419104 167994
rect 418504 131994 419104 167758
rect 418504 131758 418686 131994
rect 418922 131758 419104 131994
rect 418504 95994 419104 131758
rect 418504 95758 418686 95994
rect 418922 95758 419104 95994
rect 418504 59994 419104 95758
rect 418504 59758 418686 59994
rect 418922 59758 419104 59994
rect 418504 23994 419104 59758
rect 418504 23758 418686 23994
rect 418922 23758 419104 23994
rect 418504 -3226 419104 23758
rect 418504 -3462 418686 -3226
rect 418922 -3462 419104 -3226
rect 418504 -3546 419104 -3462
rect 418504 -3782 418686 -3546
rect 418922 -3782 419104 -3546
rect 418504 -3814 419104 -3782
rect 422204 315694 422804 338000
rect 423446 336837 423506 339630
rect 425654 337653 425714 339630
rect 425651 337652 425717 337653
rect 425651 337588 425652 337652
rect 425716 337588 425717 337652
rect 425651 337587 425717 337588
rect 423443 336836 423509 336837
rect 423443 336772 423444 336836
rect 423508 336772 423509 336836
rect 423443 336771 423509 336772
rect 422204 315458 422386 315694
rect 422622 315458 422804 315694
rect 422204 279694 422804 315458
rect 422204 279458 422386 279694
rect 422622 279458 422804 279694
rect 422204 243694 422804 279458
rect 422204 243458 422386 243694
rect 422622 243458 422804 243694
rect 422204 207694 422804 243458
rect 422204 207458 422386 207694
rect 422622 207458 422804 207694
rect 422204 171694 422804 207458
rect 422204 171458 422386 171694
rect 422622 171458 422804 171694
rect 422204 135694 422804 171458
rect 422204 135458 422386 135694
rect 422622 135458 422804 135694
rect 422204 99694 422804 135458
rect 422204 99458 422386 99694
rect 422622 99458 422804 99694
rect 422204 63694 422804 99458
rect 422204 63458 422386 63694
rect 422622 63458 422804 63694
rect 422204 27694 422804 63458
rect 422204 27458 422386 27694
rect 422622 27458 422804 27694
rect 422204 -5146 422804 27458
rect 422204 -5382 422386 -5146
rect 422622 -5382 422804 -5146
rect 422204 -5466 422804 -5382
rect 422204 -5702 422386 -5466
rect 422622 -5702 422804 -5466
rect 422204 -5734 422804 -5702
rect 425904 319394 426504 338000
rect 428598 337653 428658 339630
rect 430990 339630 431052 339690
rect 433440 339690 433500 340000
rect 435888 339690 435948 340000
rect 438472 339690 438532 340000
rect 433440 339630 433626 339690
rect 430990 337653 431050 339630
rect 428595 337652 428661 337653
rect 428595 337588 428596 337652
rect 428660 337588 428661 337652
rect 428595 337587 428661 337588
rect 430987 337652 431053 337653
rect 430987 337588 430988 337652
rect 431052 337588 431053 337652
rect 430987 337587 431053 337588
rect 425904 319158 426086 319394
rect 426322 319158 426504 319394
rect 425904 283394 426504 319158
rect 425904 283158 426086 283394
rect 426322 283158 426504 283394
rect 425904 247394 426504 283158
rect 425904 247158 426086 247394
rect 426322 247158 426504 247394
rect 425904 211394 426504 247158
rect 425904 211158 426086 211394
rect 426322 211158 426504 211394
rect 425904 175394 426504 211158
rect 425904 175158 426086 175394
rect 426322 175158 426504 175394
rect 425904 139394 426504 175158
rect 425904 139158 426086 139394
rect 426322 139158 426504 139394
rect 425904 103394 426504 139158
rect 425904 103158 426086 103394
rect 426322 103158 426504 103394
rect 425904 67394 426504 103158
rect 425904 67158 426086 67394
rect 426322 67158 426504 67394
rect 425904 31394 426504 67158
rect 425904 31158 426086 31394
rect 426322 31158 426504 31394
rect 407904 -6342 408086 -6106
rect 408322 -6342 408504 -6106
rect 407904 -6426 408504 -6342
rect 407904 -6662 408086 -6426
rect 408322 -6662 408504 -6426
rect 407904 -7654 408504 -6662
rect 425904 -7066 426504 31158
rect 432804 326294 433404 338000
rect 433566 337653 433626 339630
rect 435774 339630 435948 339690
rect 438350 339630 438532 339690
rect 440920 339690 440980 340000
rect 443368 339690 443428 340000
rect 445952 339690 446012 340000
rect 440920 339630 440986 339690
rect 433563 337652 433629 337653
rect 433563 337588 433564 337652
rect 433628 337588 433629 337652
rect 433563 337587 433629 337588
rect 435774 337109 435834 339630
rect 435771 337108 435837 337109
rect 435771 337044 435772 337108
rect 435836 337044 435837 337108
rect 435771 337043 435837 337044
rect 432804 326058 432986 326294
rect 433222 326058 433404 326294
rect 432804 290294 433404 326058
rect 432804 290058 432986 290294
rect 433222 290058 433404 290294
rect 432804 254294 433404 290058
rect 432804 254058 432986 254294
rect 433222 254058 433404 254294
rect 432804 218294 433404 254058
rect 432804 218058 432986 218294
rect 433222 218058 433404 218294
rect 432804 182294 433404 218058
rect 432804 182058 432986 182294
rect 433222 182058 433404 182294
rect 432804 146294 433404 182058
rect 432804 146058 432986 146294
rect 433222 146058 433404 146294
rect 432804 110294 433404 146058
rect 432804 110058 432986 110294
rect 433222 110058 433404 110294
rect 432804 74294 433404 110058
rect 432804 74058 432986 74294
rect 433222 74058 433404 74294
rect 432804 38294 433404 74058
rect 432804 38058 432986 38294
rect 433222 38058 433404 38294
rect 432804 2294 433404 38058
rect 432804 2058 432986 2294
rect 433222 2058 433404 2294
rect 432804 -346 433404 2058
rect 432804 -582 432986 -346
rect 433222 -582 433404 -346
rect 432804 -666 433404 -582
rect 432804 -902 432986 -666
rect 433222 -902 433404 -666
rect 432804 -1894 433404 -902
rect 436504 329994 437104 338000
rect 438350 337109 438410 339630
rect 438347 337108 438413 337109
rect 438347 337044 438348 337108
rect 438412 337044 438413 337108
rect 438347 337043 438413 337044
rect 436504 329758 436686 329994
rect 436922 329758 437104 329994
rect 436504 293994 437104 329758
rect 436504 293758 436686 293994
rect 436922 293758 437104 293994
rect 436504 257994 437104 293758
rect 436504 257758 436686 257994
rect 436922 257758 437104 257994
rect 436504 221994 437104 257758
rect 436504 221758 436686 221994
rect 436922 221758 437104 221994
rect 436504 185994 437104 221758
rect 436504 185758 436686 185994
rect 436922 185758 437104 185994
rect 436504 149994 437104 185758
rect 436504 149758 436686 149994
rect 436922 149758 437104 149994
rect 436504 113994 437104 149758
rect 436504 113758 436686 113994
rect 436922 113758 437104 113994
rect 436504 77994 437104 113758
rect 436504 77758 436686 77994
rect 436922 77758 437104 77994
rect 436504 41994 437104 77758
rect 436504 41758 436686 41994
rect 436922 41758 437104 41994
rect 436504 5994 437104 41758
rect 436504 5758 436686 5994
rect 436922 5758 437104 5994
rect 436504 -2266 437104 5758
rect 436504 -2502 436686 -2266
rect 436922 -2502 437104 -2266
rect 436504 -2586 437104 -2502
rect 436504 -2822 436686 -2586
rect 436922 -2822 437104 -2586
rect 436504 -3814 437104 -2822
rect 440204 333694 440804 338000
rect 440926 337653 440986 339630
rect 443318 339630 443428 339690
rect 445894 339630 446012 339690
rect 443318 337653 443378 339630
rect 440923 337652 440989 337653
rect 440923 337588 440924 337652
rect 440988 337588 440989 337652
rect 440923 337587 440989 337588
rect 443315 337652 443381 337653
rect 443315 337588 443316 337652
rect 443380 337588 443381 337652
rect 443315 337587 443381 337588
rect 440204 333458 440386 333694
rect 440622 333458 440804 333694
rect 440204 297694 440804 333458
rect 440204 297458 440386 297694
rect 440622 297458 440804 297694
rect 440204 261694 440804 297458
rect 440204 261458 440386 261694
rect 440622 261458 440804 261694
rect 440204 225694 440804 261458
rect 440204 225458 440386 225694
rect 440622 225458 440804 225694
rect 440204 189694 440804 225458
rect 440204 189458 440386 189694
rect 440622 189458 440804 189694
rect 440204 153694 440804 189458
rect 440204 153458 440386 153694
rect 440622 153458 440804 153694
rect 440204 117694 440804 153458
rect 440204 117458 440386 117694
rect 440622 117458 440804 117694
rect 440204 81694 440804 117458
rect 440204 81458 440386 81694
rect 440622 81458 440804 81694
rect 440204 45694 440804 81458
rect 440204 45458 440386 45694
rect 440622 45458 440804 45694
rect 440204 9694 440804 45458
rect 440204 9458 440386 9694
rect 440622 9458 440804 9694
rect 440204 -4186 440804 9458
rect 440204 -4422 440386 -4186
rect 440622 -4422 440804 -4186
rect 440204 -4506 440804 -4422
rect 440204 -4742 440386 -4506
rect 440622 -4742 440804 -4506
rect 440204 -5734 440804 -4742
rect 443904 337394 444504 338000
rect 443904 337158 444086 337394
rect 444322 337158 444504 337394
rect 445894 337245 445954 339630
rect 445891 337244 445957 337245
rect 445891 337180 445892 337244
rect 445956 337180 445957 337244
rect 445891 337179 445957 337180
rect 443904 301394 444504 337158
rect 443904 301158 444086 301394
rect 444322 301158 444504 301394
rect 443904 265394 444504 301158
rect 443904 265158 444086 265394
rect 444322 265158 444504 265394
rect 443904 229394 444504 265158
rect 443904 229158 444086 229394
rect 444322 229158 444504 229394
rect 443904 193394 444504 229158
rect 443904 193158 444086 193394
rect 444322 193158 444504 193394
rect 443904 157394 444504 193158
rect 443904 157158 444086 157394
rect 444322 157158 444504 157394
rect 443904 121394 444504 157158
rect 443904 121158 444086 121394
rect 444322 121158 444504 121394
rect 443904 85394 444504 121158
rect 443904 85158 444086 85394
rect 444322 85158 444504 85394
rect 443904 49394 444504 85158
rect 443904 49158 444086 49394
rect 444322 49158 444504 49394
rect 443904 13394 444504 49158
rect 443904 13158 444086 13394
rect 444322 13158 444504 13394
rect 425904 -7302 426086 -7066
rect 426322 -7302 426504 -7066
rect 425904 -7386 426504 -7302
rect 425904 -7622 426086 -7386
rect 426322 -7622 426504 -7386
rect 425904 -7654 426504 -7622
rect 443904 -6106 444504 13158
rect 450804 308294 451404 338000
rect 450804 308058 450986 308294
rect 451222 308058 451404 308294
rect 450804 272294 451404 308058
rect 450804 272058 450986 272294
rect 451222 272058 451404 272294
rect 450804 236294 451404 272058
rect 450804 236058 450986 236294
rect 451222 236058 451404 236294
rect 450804 200294 451404 236058
rect 450804 200058 450986 200294
rect 451222 200058 451404 200294
rect 450804 164294 451404 200058
rect 450804 164058 450986 164294
rect 451222 164058 451404 164294
rect 450804 128294 451404 164058
rect 450804 128058 450986 128294
rect 451222 128058 451404 128294
rect 450804 92294 451404 128058
rect 450804 92058 450986 92294
rect 451222 92058 451404 92294
rect 450804 56294 451404 92058
rect 450804 56058 450986 56294
rect 451222 56058 451404 56294
rect 450804 20294 451404 56058
rect 450804 20058 450986 20294
rect 451222 20058 451404 20294
rect 450804 -1306 451404 20058
rect 450804 -1542 450986 -1306
rect 451222 -1542 451404 -1306
rect 450804 -1626 451404 -1542
rect 450804 -1862 450986 -1626
rect 451222 -1862 451404 -1626
rect 450804 -1894 451404 -1862
rect 454504 311994 455104 338000
rect 454504 311758 454686 311994
rect 454922 311758 455104 311994
rect 454504 275994 455104 311758
rect 454504 275758 454686 275994
rect 454922 275758 455104 275994
rect 454504 239994 455104 275758
rect 454504 239758 454686 239994
rect 454922 239758 455104 239994
rect 454504 203994 455104 239758
rect 454504 203758 454686 203994
rect 454922 203758 455104 203994
rect 454504 167994 455104 203758
rect 454504 167758 454686 167994
rect 454922 167758 455104 167994
rect 454504 131994 455104 167758
rect 454504 131758 454686 131994
rect 454922 131758 455104 131994
rect 454504 95994 455104 131758
rect 454504 95758 454686 95994
rect 454922 95758 455104 95994
rect 454504 59994 455104 95758
rect 454504 59758 454686 59994
rect 454922 59758 455104 59994
rect 454504 23994 455104 59758
rect 454504 23758 454686 23994
rect 454922 23758 455104 23994
rect 454504 -3226 455104 23758
rect 454504 -3462 454686 -3226
rect 454922 -3462 455104 -3226
rect 454504 -3546 455104 -3462
rect 454504 -3782 454686 -3546
rect 454922 -3782 455104 -3546
rect 454504 -3814 455104 -3782
rect 458204 315694 458804 338000
rect 458204 315458 458386 315694
rect 458622 315458 458804 315694
rect 458204 279694 458804 315458
rect 458204 279458 458386 279694
rect 458622 279458 458804 279694
rect 458204 243694 458804 279458
rect 458204 243458 458386 243694
rect 458622 243458 458804 243694
rect 458204 207694 458804 243458
rect 458204 207458 458386 207694
rect 458622 207458 458804 207694
rect 458204 171694 458804 207458
rect 458204 171458 458386 171694
rect 458622 171458 458804 171694
rect 458204 135694 458804 171458
rect 458204 135458 458386 135694
rect 458622 135458 458804 135694
rect 458204 99694 458804 135458
rect 458204 99458 458386 99694
rect 458622 99458 458804 99694
rect 458204 63694 458804 99458
rect 458204 63458 458386 63694
rect 458622 63458 458804 63694
rect 458204 27694 458804 63458
rect 458204 27458 458386 27694
rect 458622 27458 458804 27694
rect 458204 -5146 458804 27458
rect 458204 -5382 458386 -5146
rect 458622 -5382 458804 -5146
rect 458204 -5466 458804 -5382
rect 458204 -5702 458386 -5466
rect 458622 -5702 458804 -5466
rect 458204 -5734 458804 -5702
rect 461904 319394 462504 338000
rect 461904 319158 462086 319394
rect 462322 319158 462504 319394
rect 461904 283394 462504 319158
rect 461904 283158 462086 283394
rect 462322 283158 462504 283394
rect 461904 247394 462504 283158
rect 461904 247158 462086 247394
rect 462322 247158 462504 247394
rect 461904 211394 462504 247158
rect 461904 211158 462086 211394
rect 462322 211158 462504 211394
rect 461904 175394 462504 211158
rect 461904 175158 462086 175394
rect 462322 175158 462504 175394
rect 461904 139394 462504 175158
rect 461904 139158 462086 139394
rect 462322 139158 462504 139394
rect 461904 103394 462504 139158
rect 461904 103158 462086 103394
rect 462322 103158 462504 103394
rect 461904 67394 462504 103158
rect 461904 67158 462086 67394
rect 462322 67158 462504 67394
rect 461904 31394 462504 67158
rect 461904 31158 462086 31394
rect 462322 31158 462504 31394
rect 443904 -6342 444086 -6106
rect 444322 -6342 444504 -6106
rect 443904 -6426 444504 -6342
rect 443904 -6662 444086 -6426
rect 444322 -6662 444504 -6426
rect 443904 -7654 444504 -6662
rect 461904 -7066 462504 31158
rect 468804 326294 469404 338000
rect 468804 326058 468986 326294
rect 469222 326058 469404 326294
rect 468804 290294 469404 326058
rect 468804 290058 468986 290294
rect 469222 290058 469404 290294
rect 468804 254294 469404 290058
rect 468804 254058 468986 254294
rect 469222 254058 469404 254294
rect 468804 218294 469404 254058
rect 468804 218058 468986 218294
rect 469222 218058 469404 218294
rect 468804 182294 469404 218058
rect 468804 182058 468986 182294
rect 469222 182058 469404 182294
rect 468804 146294 469404 182058
rect 468804 146058 468986 146294
rect 469222 146058 469404 146294
rect 468804 110294 469404 146058
rect 468804 110058 468986 110294
rect 469222 110058 469404 110294
rect 468804 74294 469404 110058
rect 468804 74058 468986 74294
rect 469222 74058 469404 74294
rect 468804 38294 469404 74058
rect 468804 38058 468986 38294
rect 469222 38058 469404 38294
rect 468804 2294 469404 38058
rect 468804 2058 468986 2294
rect 469222 2058 469404 2294
rect 468804 -346 469404 2058
rect 468804 -582 468986 -346
rect 469222 -582 469404 -346
rect 468804 -666 469404 -582
rect 468804 -902 468986 -666
rect 469222 -902 469404 -666
rect 468804 -1894 469404 -902
rect 472504 329994 473104 338000
rect 472504 329758 472686 329994
rect 472922 329758 473104 329994
rect 472504 293994 473104 329758
rect 472504 293758 472686 293994
rect 472922 293758 473104 293994
rect 472504 257994 473104 293758
rect 472504 257758 472686 257994
rect 472922 257758 473104 257994
rect 472504 221994 473104 257758
rect 472504 221758 472686 221994
rect 472922 221758 473104 221994
rect 472504 185994 473104 221758
rect 472504 185758 472686 185994
rect 472922 185758 473104 185994
rect 472504 149994 473104 185758
rect 472504 149758 472686 149994
rect 472922 149758 473104 149994
rect 472504 113994 473104 149758
rect 472504 113758 472686 113994
rect 472922 113758 473104 113994
rect 472504 77994 473104 113758
rect 472504 77758 472686 77994
rect 472922 77758 473104 77994
rect 472504 41994 473104 77758
rect 472504 41758 472686 41994
rect 472922 41758 473104 41994
rect 472504 5994 473104 41758
rect 472504 5758 472686 5994
rect 472922 5758 473104 5994
rect 472504 -2266 473104 5758
rect 472504 -2502 472686 -2266
rect 472922 -2502 473104 -2266
rect 472504 -2586 473104 -2502
rect 472504 -2822 472686 -2586
rect 472922 -2822 473104 -2586
rect 472504 -3814 473104 -2822
rect 476204 333694 476804 338000
rect 476204 333458 476386 333694
rect 476622 333458 476804 333694
rect 476204 297694 476804 333458
rect 476204 297458 476386 297694
rect 476622 297458 476804 297694
rect 476204 261694 476804 297458
rect 476204 261458 476386 261694
rect 476622 261458 476804 261694
rect 476204 225694 476804 261458
rect 476204 225458 476386 225694
rect 476622 225458 476804 225694
rect 476204 189694 476804 225458
rect 476204 189458 476386 189694
rect 476622 189458 476804 189694
rect 476204 153694 476804 189458
rect 476204 153458 476386 153694
rect 476622 153458 476804 153694
rect 476204 117694 476804 153458
rect 476204 117458 476386 117694
rect 476622 117458 476804 117694
rect 476204 81694 476804 117458
rect 476204 81458 476386 81694
rect 476622 81458 476804 81694
rect 476204 45694 476804 81458
rect 476204 45458 476386 45694
rect 476622 45458 476804 45694
rect 476204 9694 476804 45458
rect 476204 9458 476386 9694
rect 476622 9458 476804 9694
rect 476204 -4186 476804 9458
rect 476204 -4422 476386 -4186
rect 476622 -4422 476804 -4186
rect 476204 -4506 476804 -4422
rect 476204 -4742 476386 -4506
rect 476622 -4742 476804 -4506
rect 476204 -5734 476804 -4742
rect 479904 337394 480504 373158
rect 479904 337158 480086 337394
rect 480322 337158 480504 337394
rect 479904 301394 480504 337158
rect 479904 301158 480086 301394
rect 480322 301158 480504 301394
rect 479904 265394 480504 301158
rect 479904 265158 480086 265394
rect 480322 265158 480504 265394
rect 479904 229394 480504 265158
rect 479904 229158 480086 229394
rect 480322 229158 480504 229394
rect 479904 193394 480504 229158
rect 479904 193158 480086 193394
rect 480322 193158 480504 193394
rect 479904 157394 480504 193158
rect 479904 157158 480086 157394
rect 480322 157158 480504 157394
rect 479904 121394 480504 157158
rect 479904 121158 480086 121394
rect 480322 121158 480504 121394
rect 479904 85394 480504 121158
rect 479904 85158 480086 85394
rect 480322 85158 480504 85394
rect 479904 49394 480504 85158
rect 479904 49158 480086 49394
rect 480322 49158 480504 49394
rect 479904 13394 480504 49158
rect 479904 13158 480086 13394
rect 480322 13158 480504 13394
rect 461904 -7302 462086 -7066
rect 462322 -7302 462504 -7066
rect 461904 -7386 462504 -7302
rect 461904 -7622 462086 -7386
rect 462322 -7622 462504 -7386
rect 461904 -7654 462504 -7622
rect 479904 -6106 480504 13158
rect 486804 705798 487404 705830
rect 486804 705562 486986 705798
rect 487222 705562 487404 705798
rect 486804 705478 487404 705562
rect 486804 705242 486986 705478
rect 487222 705242 487404 705478
rect 486804 668294 487404 705242
rect 486804 668058 486986 668294
rect 487222 668058 487404 668294
rect 486804 632294 487404 668058
rect 486804 632058 486986 632294
rect 487222 632058 487404 632294
rect 486804 596294 487404 632058
rect 486804 596058 486986 596294
rect 487222 596058 487404 596294
rect 486804 560294 487404 596058
rect 486804 560058 486986 560294
rect 487222 560058 487404 560294
rect 486804 524294 487404 560058
rect 486804 524058 486986 524294
rect 487222 524058 487404 524294
rect 486804 488294 487404 524058
rect 486804 488058 486986 488294
rect 487222 488058 487404 488294
rect 486804 452294 487404 488058
rect 486804 452058 486986 452294
rect 487222 452058 487404 452294
rect 486804 416294 487404 452058
rect 486804 416058 486986 416294
rect 487222 416058 487404 416294
rect 486804 380294 487404 416058
rect 486804 380058 486986 380294
rect 487222 380058 487404 380294
rect 486804 344294 487404 380058
rect 486804 344058 486986 344294
rect 487222 344058 487404 344294
rect 486804 308294 487404 344058
rect 486804 308058 486986 308294
rect 487222 308058 487404 308294
rect 486804 272294 487404 308058
rect 486804 272058 486986 272294
rect 487222 272058 487404 272294
rect 486804 236294 487404 272058
rect 486804 236058 486986 236294
rect 487222 236058 487404 236294
rect 486804 200294 487404 236058
rect 486804 200058 486986 200294
rect 487222 200058 487404 200294
rect 486804 164294 487404 200058
rect 486804 164058 486986 164294
rect 487222 164058 487404 164294
rect 486804 128294 487404 164058
rect 486804 128058 486986 128294
rect 487222 128058 487404 128294
rect 486804 92294 487404 128058
rect 486804 92058 486986 92294
rect 487222 92058 487404 92294
rect 486804 56294 487404 92058
rect 486804 56058 486986 56294
rect 487222 56058 487404 56294
rect 486804 20294 487404 56058
rect 486804 20058 486986 20294
rect 487222 20058 487404 20294
rect 486804 -1306 487404 20058
rect 486804 -1542 486986 -1306
rect 487222 -1542 487404 -1306
rect 486804 -1626 487404 -1542
rect 486804 -1862 486986 -1626
rect 487222 -1862 487404 -1626
rect 486804 -1894 487404 -1862
rect 490504 671994 491104 707162
rect 490504 671758 490686 671994
rect 490922 671758 491104 671994
rect 490504 635994 491104 671758
rect 490504 635758 490686 635994
rect 490922 635758 491104 635994
rect 490504 599994 491104 635758
rect 490504 599758 490686 599994
rect 490922 599758 491104 599994
rect 490504 563994 491104 599758
rect 490504 563758 490686 563994
rect 490922 563758 491104 563994
rect 490504 527994 491104 563758
rect 490504 527758 490686 527994
rect 490922 527758 491104 527994
rect 490504 491994 491104 527758
rect 490504 491758 490686 491994
rect 490922 491758 491104 491994
rect 490504 455994 491104 491758
rect 490504 455758 490686 455994
rect 490922 455758 491104 455994
rect 490504 419994 491104 455758
rect 490504 419758 490686 419994
rect 490922 419758 491104 419994
rect 490504 383994 491104 419758
rect 490504 383758 490686 383994
rect 490922 383758 491104 383994
rect 490504 347994 491104 383758
rect 490504 347758 490686 347994
rect 490922 347758 491104 347994
rect 490504 311994 491104 347758
rect 490504 311758 490686 311994
rect 490922 311758 491104 311994
rect 490504 275994 491104 311758
rect 490504 275758 490686 275994
rect 490922 275758 491104 275994
rect 490504 239994 491104 275758
rect 490504 239758 490686 239994
rect 490922 239758 491104 239994
rect 490504 203994 491104 239758
rect 490504 203758 490686 203994
rect 490922 203758 491104 203994
rect 490504 167994 491104 203758
rect 490504 167758 490686 167994
rect 490922 167758 491104 167994
rect 490504 131994 491104 167758
rect 490504 131758 490686 131994
rect 490922 131758 491104 131994
rect 490504 95994 491104 131758
rect 490504 95758 490686 95994
rect 490922 95758 491104 95994
rect 490504 59994 491104 95758
rect 490504 59758 490686 59994
rect 490922 59758 491104 59994
rect 490504 23994 491104 59758
rect 490504 23758 490686 23994
rect 490922 23758 491104 23994
rect 490504 -3226 491104 23758
rect 490504 -3462 490686 -3226
rect 490922 -3462 491104 -3226
rect 490504 -3546 491104 -3462
rect 490504 -3782 490686 -3546
rect 490922 -3782 491104 -3546
rect 490504 -3814 491104 -3782
rect 494204 675694 494804 709082
rect 494204 675458 494386 675694
rect 494622 675458 494804 675694
rect 494204 639694 494804 675458
rect 494204 639458 494386 639694
rect 494622 639458 494804 639694
rect 494204 603694 494804 639458
rect 494204 603458 494386 603694
rect 494622 603458 494804 603694
rect 494204 567694 494804 603458
rect 494204 567458 494386 567694
rect 494622 567458 494804 567694
rect 494204 531694 494804 567458
rect 494204 531458 494386 531694
rect 494622 531458 494804 531694
rect 494204 495694 494804 531458
rect 494204 495458 494386 495694
rect 494622 495458 494804 495694
rect 494204 459694 494804 495458
rect 494204 459458 494386 459694
rect 494622 459458 494804 459694
rect 494204 423694 494804 459458
rect 494204 423458 494386 423694
rect 494622 423458 494804 423694
rect 494204 387694 494804 423458
rect 494204 387458 494386 387694
rect 494622 387458 494804 387694
rect 494204 351694 494804 387458
rect 494204 351458 494386 351694
rect 494622 351458 494804 351694
rect 494204 315694 494804 351458
rect 494204 315458 494386 315694
rect 494622 315458 494804 315694
rect 494204 279694 494804 315458
rect 494204 279458 494386 279694
rect 494622 279458 494804 279694
rect 494204 243694 494804 279458
rect 494204 243458 494386 243694
rect 494622 243458 494804 243694
rect 494204 207694 494804 243458
rect 494204 207458 494386 207694
rect 494622 207458 494804 207694
rect 494204 171694 494804 207458
rect 494204 171458 494386 171694
rect 494622 171458 494804 171694
rect 494204 135694 494804 171458
rect 494204 135458 494386 135694
rect 494622 135458 494804 135694
rect 494204 99694 494804 135458
rect 494204 99458 494386 99694
rect 494622 99458 494804 99694
rect 494204 63694 494804 99458
rect 494204 63458 494386 63694
rect 494622 63458 494804 63694
rect 494204 27694 494804 63458
rect 494204 27458 494386 27694
rect 494622 27458 494804 27694
rect 494204 -5146 494804 27458
rect 494204 -5382 494386 -5146
rect 494622 -5382 494804 -5146
rect 494204 -5466 494804 -5382
rect 494204 -5702 494386 -5466
rect 494622 -5702 494804 -5466
rect 494204 -5734 494804 -5702
rect 497904 679394 498504 711002
rect 515904 710598 516504 711590
rect 515904 710362 516086 710598
rect 516322 710362 516504 710598
rect 515904 710278 516504 710362
rect 515904 710042 516086 710278
rect 516322 710042 516504 710278
rect 512204 708678 512804 709670
rect 512204 708442 512386 708678
rect 512622 708442 512804 708678
rect 512204 708358 512804 708442
rect 512204 708122 512386 708358
rect 512622 708122 512804 708358
rect 508504 706758 509104 707750
rect 508504 706522 508686 706758
rect 508922 706522 509104 706758
rect 508504 706438 509104 706522
rect 508504 706202 508686 706438
rect 508922 706202 509104 706438
rect 497904 679158 498086 679394
rect 498322 679158 498504 679394
rect 497904 643394 498504 679158
rect 497904 643158 498086 643394
rect 498322 643158 498504 643394
rect 497904 607394 498504 643158
rect 497904 607158 498086 607394
rect 498322 607158 498504 607394
rect 497904 571394 498504 607158
rect 497904 571158 498086 571394
rect 498322 571158 498504 571394
rect 497904 535394 498504 571158
rect 497904 535158 498086 535394
rect 498322 535158 498504 535394
rect 497904 499394 498504 535158
rect 497904 499158 498086 499394
rect 498322 499158 498504 499394
rect 497904 463394 498504 499158
rect 497904 463158 498086 463394
rect 498322 463158 498504 463394
rect 497904 427394 498504 463158
rect 497904 427158 498086 427394
rect 498322 427158 498504 427394
rect 497904 391394 498504 427158
rect 497904 391158 498086 391394
rect 498322 391158 498504 391394
rect 497904 355394 498504 391158
rect 497904 355158 498086 355394
rect 498322 355158 498504 355394
rect 497904 319394 498504 355158
rect 497904 319158 498086 319394
rect 498322 319158 498504 319394
rect 497904 283394 498504 319158
rect 497904 283158 498086 283394
rect 498322 283158 498504 283394
rect 497904 247394 498504 283158
rect 497904 247158 498086 247394
rect 498322 247158 498504 247394
rect 497904 211394 498504 247158
rect 497904 211158 498086 211394
rect 498322 211158 498504 211394
rect 497904 175394 498504 211158
rect 497904 175158 498086 175394
rect 498322 175158 498504 175394
rect 497904 139394 498504 175158
rect 497904 139158 498086 139394
rect 498322 139158 498504 139394
rect 497904 103394 498504 139158
rect 497904 103158 498086 103394
rect 498322 103158 498504 103394
rect 497904 67394 498504 103158
rect 497904 67158 498086 67394
rect 498322 67158 498504 67394
rect 497904 31394 498504 67158
rect 497904 31158 498086 31394
rect 498322 31158 498504 31394
rect 479904 -6342 480086 -6106
rect 480322 -6342 480504 -6106
rect 479904 -6426 480504 -6342
rect 479904 -6662 480086 -6426
rect 480322 -6662 480504 -6426
rect 479904 -7654 480504 -6662
rect 497904 -7066 498504 31158
rect 504804 704838 505404 705830
rect 504804 704602 504986 704838
rect 505222 704602 505404 704838
rect 504804 704518 505404 704602
rect 504804 704282 504986 704518
rect 505222 704282 505404 704518
rect 504804 686294 505404 704282
rect 504804 686058 504986 686294
rect 505222 686058 505404 686294
rect 504804 650294 505404 686058
rect 504804 650058 504986 650294
rect 505222 650058 505404 650294
rect 504804 614294 505404 650058
rect 504804 614058 504986 614294
rect 505222 614058 505404 614294
rect 504804 578294 505404 614058
rect 504804 578058 504986 578294
rect 505222 578058 505404 578294
rect 504804 542294 505404 578058
rect 504804 542058 504986 542294
rect 505222 542058 505404 542294
rect 504804 506294 505404 542058
rect 504804 506058 504986 506294
rect 505222 506058 505404 506294
rect 504804 470294 505404 506058
rect 504804 470058 504986 470294
rect 505222 470058 505404 470294
rect 504804 434294 505404 470058
rect 504804 434058 504986 434294
rect 505222 434058 505404 434294
rect 504804 398294 505404 434058
rect 504804 398058 504986 398294
rect 505222 398058 505404 398294
rect 504804 362294 505404 398058
rect 504804 362058 504986 362294
rect 505222 362058 505404 362294
rect 504804 326294 505404 362058
rect 504804 326058 504986 326294
rect 505222 326058 505404 326294
rect 504804 290294 505404 326058
rect 504804 290058 504986 290294
rect 505222 290058 505404 290294
rect 504804 254294 505404 290058
rect 504804 254058 504986 254294
rect 505222 254058 505404 254294
rect 504804 218294 505404 254058
rect 504804 218058 504986 218294
rect 505222 218058 505404 218294
rect 504804 182294 505404 218058
rect 504804 182058 504986 182294
rect 505222 182058 505404 182294
rect 504804 146294 505404 182058
rect 504804 146058 504986 146294
rect 505222 146058 505404 146294
rect 504804 110294 505404 146058
rect 504804 110058 504986 110294
rect 505222 110058 505404 110294
rect 504804 74294 505404 110058
rect 504804 74058 504986 74294
rect 505222 74058 505404 74294
rect 504804 38294 505404 74058
rect 504804 38058 504986 38294
rect 505222 38058 505404 38294
rect 504804 2294 505404 38058
rect 504804 2058 504986 2294
rect 505222 2058 505404 2294
rect 504804 -346 505404 2058
rect 504804 -582 504986 -346
rect 505222 -582 505404 -346
rect 504804 -666 505404 -582
rect 504804 -902 504986 -666
rect 505222 -902 505404 -666
rect 504804 -1894 505404 -902
rect 508504 689994 509104 706202
rect 508504 689758 508686 689994
rect 508922 689758 509104 689994
rect 508504 653994 509104 689758
rect 508504 653758 508686 653994
rect 508922 653758 509104 653994
rect 508504 617994 509104 653758
rect 508504 617758 508686 617994
rect 508922 617758 509104 617994
rect 508504 581994 509104 617758
rect 508504 581758 508686 581994
rect 508922 581758 509104 581994
rect 508504 545994 509104 581758
rect 508504 545758 508686 545994
rect 508922 545758 509104 545994
rect 508504 509994 509104 545758
rect 508504 509758 508686 509994
rect 508922 509758 509104 509994
rect 508504 473994 509104 509758
rect 508504 473758 508686 473994
rect 508922 473758 509104 473994
rect 508504 437994 509104 473758
rect 508504 437758 508686 437994
rect 508922 437758 509104 437994
rect 508504 401994 509104 437758
rect 508504 401758 508686 401994
rect 508922 401758 509104 401994
rect 508504 365994 509104 401758
rect 508504 365758 508686 365994
rect 508922 365758 509104 365994
rect 508504 329994 509104 365758
rect 508504 329758 508686 329994
rect 508922 329758 509104 329994
rect 508504 293994 509104 329758
rect 508504 293758 508686 293994
rect 508922 293758 509104 293994
rect 508504 257994 509104 293758
rect 508504 257758 508686 257994
rect 508922 257758 509104 257994
rect 508504 221994 509104 257758
rect 508504 221758 508686 221994
rect 508922 221758 509104 221994
rect 508504 185994 509104 221758
rect 508504 185758 508686 185994
rect 508922 185758 509104 185994
rect 508504 149994 509104 185758
rect 508504 149758 508686 149994
rect 508922 149758 509104 149994
rect 508504 113994 509104 149758
rect 508504 113758 508686 113994
rect 508922 113758 509104 113994
rect 508504 77994 509104 113758
rect 508504 77758 508686 77994
rect 508922 77758 509104 77994
rect 508504 41994 509104 77758
rect 508504 41758 508686 41994
rect 508922 41758 509104 41994
rect 508504 5994 509104 41758
rect 508504 5758 508686 5994
rect 508922 5758 509104 5994
rect 508504 -2266 509104 5758
rect 508504 -2502 508686 -2266
rect 508922 -2502 509104 -2266
rect 508504 -2586 509104 -2502
rect 508504 -2822 508686 -2586
rect 508922 -2822 509104 -2586
rect 508504 -3814 509104 -2822
rect 512204 693694 512804 708122
rect 512204 693458 512386 693694
rect 512622 693458 512804 693694
rect 512204 657694 512804 693458
rect 512204 657458 512386 657694
rect 512622 657458 512804 657694
rect 512204 621694 512804 657458
rect 512204 621458 512386 621694
rect 512622 621458 512804 621694
rect 512204 585694 512804 621458
rect 512204 585458 512386 585694
rect 512622 585458 512804 585694
rect 512204 549694 512804 585458
rect 512204 549458 512386 549694
rect 512622 549458 512804 549694
rect 512204 513694 512804 549458
rect 512204 513458 512386 513694
rect 512622 513458 512804 513694
rect 512204 477694 512804 513458
rect 512204 477458 512386 477694
rect 512622 477458 512804 477694
rect 512204 441694 512804 477458
rect 512204 441458 512386 441694
rect 512622 441458 512804 441694
rect 512204 405694 512804 441458
rect 512204 405458 512386 405694
rect 512622 405458 512804 405694
rect 512204 369694 512804 405458
rect 512204 369458 512386 369694
rect 512622 369458 512804 369694
rect 512204 333694 512804 369458
rect 512204 333458 512386 333694
rect 512622 333458 512804 333694
rect 512204 297694 512804 333458
rect 512204 297458 512386 297694
rect 512622 297458 512804 297694
rect 512204 261694 512804 297458
rect 512204 261458 512386 261694
rect 512622 261458 512804 261694
rect 512204 225694 512804 261458
rect 512204 225458 512386 225694
rect 512622 225458 512804 225694
rect 512204 189694 512804 225458
rect 512204 189458 512386 189694
rect 512622 189458 512804 189694
rect 512204 153694 512804 189458
rect 512204 153458 512386 153694
rect 512622 153458 512804 153694
rect 512204 117694 512804 153458
rect 512204 117458 512386 117694
rect 512622 117458 512804 117694
rect 512204 81694 512804 117458
rect 512204 81458 512386 81694
rect 512622 81458 512804 81694
rect 512204 45694 512804 81458
rect 512204 45458 512386 45694
rect 512622 45458 512804 45694
rect 512204 9694 512804 45458
rect 512204 9458 512386 9694
rect 512622 9458 512804 9694
rect 512204 -4186 512804 9458
rect 512204 -4422 512386 -4186
rect 512622 -4422 512804 -4186
rect 512204 -4506 512804 -4422
rect 512204 -4742 512386 -4506
rect 512622 -4742 512804 -4506
rect 512204 -5734 512804 -4742
rect 515904 697394 516504 710042
rect 533904 711558 534504 711590
rect 533904 711322 534086 711558
rect 534322 711322 534504 711558
rect 533904 711238 534504 711322
rect 533904 711002 534086 711238
rect 534322 711002 534504 711238
rect 530204 709638 530804 709670
rect 530204 709402 530386 709638
rect 530622 709402 530804 709638
rect 530204 709318 530804 709402
rect 530204 709082 530386 709318
rect 530622 709082 530804 709318
rect 526504 707718 527104 707750
rect 526504 707482 526686 707718
rect 526922 707482 527104 707718
rect 526504 707398 527104 707482
rect 526504 707162 526686 707398
rect 526922 707162 527104 707398
rect 515904 697158 516086 697394
rect 516322 697158 516504 697394
rect 515904 661394 516504 697158
rect 515904 661158 516086 661394
rect 516322 661158 516504 661394
rect 515904 625394 516504 661158
rect 515904 625158 516086 625394
rect 516322 625158 516504 625394
rect 515904 589394 516504 625158
rect 515904 589158 516086 589394
rect 516322 589158 516504 589394
rect 515904 553394 516504 589158
rect 515904 553158 516086 553394
rect 516322 553158 516504 553394
rect 515904 517394 516504 553158
rect 515904 517158 516086 517394
rect 516322 517158 516504 517394
rect 515904 481394 516504 517158
rect 515904 481158 516086 481394
rect 516322 481158 516504 481394
rect 515904 445394 516504 481158
rect 515904 445158 516086 445394
rect 516322 445158 516504 445394
rect 515904 409394 516504 445158
rect 515904 409158 516086 409394
rect 516322 409158 516504 409394
rect 515904 373394 516504 409158
rect 515904 373158 516086 373394
rect 516322 373158 516504 373394
rect 515904 337394 516504 373158
rect 515904 337158 516086 337394
rect 516322 337158 516504 337394
rect 515904 301394 516504 337158
rect 515904 301158 516086 301394
rect 516322 301158 516504 301394
rect 515904 265394 516504 301158
rect 515904 265158 516086 265394
rect 516322 265158 516504 265394
rect 515904 229394 516504 265158
rect 515904 229158 516086 229394
rect 516322 229158 516504 229394
rect 515904 193394 516504 229158
rect 515904 193158 516086 193394
rect 516322 193158 516504 193394
rect 515904 157394 516504 193158
rect 515904 157158 516086 157394
rect 516322 157158 516504 157394
rect 515904 121394 516504 157158
rect 515904 121158 516086 121394
rect 516322 121158 516504 121394
rect 515904 85394 516504 121158
rect 515904 85158 516086 85394
rect 516322 85158 516504 85394
rect 515904 49394 516504 85158
rect 515904 49158 516086 49394
rect 516322 49158 516504 49394
rect 515904 13394 516504 49158
rect 515904 13158 516086 13394
rect 516322 13158 516504 13394
rect 497904 -7302 498086 -7066
rect 498322 -7302 498504 -7066
rect 497904 -7386 498504 -7302
rect 497904 -7622 498086 -7386
rect 498322 -7622 498504 -7386
rect 497904 -7654 498504 -7622
rect 515904 -6106 516504 13158
rect 522804 705798 523404 705830
rect 522804 705562 522986 705798
rect 523222 705562 523404 705798
rect 522804 705478 523404 705562
rect 522804 705242 522986 705478
rect 523222 705242 523404 705478
rect 522804 668294 523404 705242
rect 522804 668058 522986 668294
rect 523222 668058 523404 668294
rect 522804 632294 523404 668058
rect 522804 632058 522986 632294
rect 523222 632058 523404 632294
rect 522804 596294 523404 632058
rect 522804 596058 522986 596294
rect 523222 596058 523404 596294
rect 522804 560294 523404 596058
rect 522804 560058 522986 560294
rect 523222 560058 523404 560294
rect 522804 524294 523404 560058
rect 522804 524058 522986 524294
rect 523222 524058 523404 524294
rect 522804 488294 523404 524058
rect 522804 488058 522986 488294
rect 523222 488058 523404 488294
rect 522804 452294 523404 488058
rect 522804 452058 522986 452294
rect 523222 452058 523404 452294
rect 522804 416294 523404 452058
rect 522804 416058 522986 416294
rect 523222 416058 523404 416294
rect 522804 380294 523404 416058
rect 522804 380058 522986 380294
rect 523222 380058 523404 380294
rect 522804 344294 523404 380058
rect 522804 344058 522986 344294
rect 523222 344058 523404 344294
rect 522804 308294 523404 344058
rect 522804 308058 522986 308294
rect 523222 308058 523404 308294
rect 522804 272294 523404 308058
rect 522804 272058 522986 272294
rect 523222 272058 523404 272294
rect 522804 236294 523404 272058
rect 522804 236058 522986 236294
rect 523222 236058 523404 236294
rect 522804 200294 523404 236058
rect 522804 200058 522986 200294
rect 523222 200058 523404 200294
rect 522804 164294 523404 200058
rect 522804 164058 522986 164294
rect 523222 164058 523404 164294
rect 522804 128294 523404 164058
rect 522804 128058 522986 128294
rect 523222 128058 523404 128294
rect 522804 92294 523404 128058
rect 522804 92058 522986 92294
rect 523222 92058 523404 92294
rect 522804 56294 523404 92058
rect 522804 56058 522986 56294
rect 523222 56058 523404 56294
rect 522804 20294 523404 56058
rect 522804 20058 522986 20294
rect 523222 20058 523404 20294
rect 522804 -1306 523404 20058
rect 522804 -1542 522986 -1306
rect 523222 -1542 523404 -1306
rect 522804 -1626 523404 -1542
rect 522804 -1862 522986 -1626
rect 523222 -1862 523404 -1626
rect 522804 -1894 523404 -1862
rect 526504 671994 527104 707162
rect 526504 671758 526686 671994
rect 526922 671758 527104 671994
rect 526504 635994 527104 671758
rect 526504 635758 526686 635994
rect 526922 635758 527104 635994
rect 526504 599994 527104 635758
rect 526504 599758 526686 599994
rect 526922 599758 527104 599994
rect 526504 563994 527104 599758
rect 526504 563758 526686 563994
rect 526922 563758 527104 563994
rect 526504 527994 527104 563758
rect 526504 527758 526686 527994
rect 526922 527758 527104 527994
rect 526504 491994 527104 527758
rect 526504 491758 526686 491994
rect 526922 491758 527104 491994
rect 526504 455994 527104 491758
rect 526504 455758 526686 455994
rect 526922 455758 527104 455994
rect 526504 419994 527104 455758
rect 526504 419758 526686 419994
rect 526922 419758 527104 419994
rect 526504 383994 527104 419758
rect 526504 383758 526686 383994
rect 526922 383758 527104 383994
rect 526504 347994 527104 383758
rect 526504 347758 526686 347994
rect 526922 347758 527104 347994
rect 526504 311994 527104 347758
rect 526504 311758 526686 311994
rect 526922 311758 527104 311994
rect 526504 275994 527104 311758
rect 526504 275758 526686 275994
rect 526922 275758 527104 275994
rect 526504 239994 527104 275758
rect 526504 239758 526686 239994
rect 526922 239758 527104 239994
rect 526504 203994 527104 239758
rect 526504 203758 526686 203994
rect 526922 203758 527104 203994
rect 526504 167994 527104 203758
rect 526504 167758 526686 167994
rect 526922 167758 527104 167994
rect 526504 131994 527104 167758
rect 526504 131758 526686 131994
rect 526922 131758 527104 131994
rect 526504 95994 527104 131758
rect 526504 95758 526686 95994
rect 526922 95758 527104 95994
rect 526504 59994 527104 95758
rect 526504 59758 526686 59994
rect 526922 59758 527104 59994
rect 526504 23994 527104 59758
rect 526504 23758 526686 23994
rect 526922 23758 527104 23994
rect 526504 -3226 527104 23758
rect 526504 -3462 526686 -3226
rect 526922 -3462 527104 -3226
rect 526504 -3546 527104 -3462
rect 526504 -3782 526686 -3546
rect 526922 -3782 527104 -3546
rect 526504 -3814 527104 -3782
rect 530204 675694 530804 709082
rect 530204 675458 530386 675694
rect 530622 675458 530804 675694
rect 530204 639694 530804 675458
rect 530204 639458 530386 639694
rect 530622 639458 530804 639694
rect 530204 603694 530804 639458
rect 530204 603458 530386 603694
rect 530622 603458 530804 603694
rect 530204 567694 530804 603458
rect 530204 567458 530386 567694
rect 530622 567458 530804 567694
rect 530204 531694 530804 567458
rect 530204 531458 530386 531694
rect 530622 531458 530804 531694
rect 530204 495694 530804 531458
rect 530204 495458 530386 495694
rect 530622 495458 530804 495694
rect 530204 459694 530804 495458
rect 530204 459458 530386 459694
rect 530622 459458 530804 459694
rect 530204 423694 530804 459458
rect 530204 423458 530386 423694
rect 530622 423458 530804 423694
rect 530204 387694 530804 423458
rect 530204 387458 530386 387694
rect 530622 387458 530804 387694
rect 530204 351694 530804 387458
rect 530204 351458 530386 351694
rect 530622 351458 530804 351694
rect 530204 315694 530804 351458
rect 530204 315458 530386 315694
rect 530622 315458 530804 315694
rect 530204 279694 530804 315458
rect 530204 279458 530386 279694
rect 530622 279458 530804 279694
rect 530204 243694 530804 279458
rect 530204 243458 530386 243694
rect 530622 243458 530804 243694
rect 530204 207694 530804 243458
rect 530204 207458 530386 207694
rect 530622 207458 530804 207694
rect 530204 171694 530804 207458
rect 530204 171458 530386 171694
rect 530622 171458 530804 171694
rect 530204 135694 530804 171458
rect 530204 135458 530386 135694
rect 530622 135458 530804 135694
rect 530204 99694 530804 135458
rect 530204 99458 530386 99694
rect 530622 99458 530804 99694
rect 530204 63694 530804 99458
rect 530204 63458 530386 63694
rect 530622 63458 530804 63694
rect 530204 27694 530804 63458
rect 530204 27458 530386 27694
rect 530622 27458 530804 27694
rect 530204 -5146 530804 27458
rect 530204 -5382 530386 -5146
rect 530622 -5382 530804 -5146
rect 530204 -5466 530804 -5382
rect 530204 -5702 530386 -5466
rect 530622 -5702 530804 -5466
rect 530204 -5734 530804 -5702
rect 533904 679394 534504 711002
rect 551904 710598 552504 711590
rect 551904 710362 552086 710598
rect 552322 710362 552504 710598
rect 551904 710278 552504 710362
rect 551904 710042 552086 710278
rect 552322 710042 552504 710278
rect 548204 708678 548804 709670
rect 548204 708442 548386 708678
rect 548622 708442 548804 708678
rect 548204 708358 548804 708442
rect 548204 708122 548386 708358
rect 548622 708122 548804 708358
rect 544504 706758 545104 707750
rect 544504 706522 544686 706758
rect 544922 706522 545104 706758
rect 544504 706438 545104 706522
rect 544504 706202 544686 706438
rect 544922 706202 545104 706438
rect 533904 679158 534086 679394
rect 534322 679158 534504 679394
rect 533904 643394 534504 679158
rect 533904 643158 534086 643394
rect 534322 643158 534504 643394
rect 533904 607394 534504 643158
rect 533904 607158 534086 607394
rect 534322 607158 534504 607394
rect 533904 571394 534504 607158
rect 533904 571158 534086 571394
rect 534322 571158 534504 571394
rect 533904 535394 534504 571158
rect 533904 535158 534086 535394
rect 534322 535158 534504 535394
rect 533904 499394 534504 535158
rect 533904 499158 534086 499394
rect 534322 499158 534504 499394
rect 533904 463394 534504 499158
rect 533904 463158 534086 463394
rect 534322 463158 534504 463394
rect 533904 427394 534504 463158
rect 533904 427158 534086 427394
rect 534322 427158 534504 427394
rect 533904 391394 534504 427158
rect 533904 391158 534086 391394
rect 534322 391158 534504 391394
rect 533904 355394 534504 391158
rect 533904 355158 534086 355394
rect 534322 355158 534504 355394
rect 533904 319394 534504 355158
rect 533904 319158 534086 319394
rect 534322 319158 534504 319394
rect 533904 283394 534504 319158
rect 533904 283158 534086 283394
rect 534322 283158 534504 283394
rect 533904 247394 534504 283158
rect 533904 247158 534086 247394
rect 534322 247158 534504 247394
rect 533904 211394 534504 247158
rect 533904 211158 534086 211394
rect 534322 211158 534504 211394
rect 533904 175394 534504 211158
rect 533904 175158 534086 175394
rect 534322 175158 534504 175394
rect 533904 139394 534504 175158
rect 533904 139158 534086 139394
rect 534322 139158 534504 139394
rect 533904 103394 534504 139158
rect 533904 103158 534086 103394
rect 534322 103158 534504 103394
rect 533904 67394 534504 103158
rect 533904 67158 534086 67394
rect 534322 67158 534504 67394
rect 533904 31394 534504 67158
rect 533904 31158 534086 31394
rect 534322 31158 534504 31394
rect 515904 -6342 516086 -6106
rect 516322 -6342 516504 -6106
rect 515904 -6426 516504 -6342
rect 515904 -6662 516086 -6426
rect 516322 -6662 516504 -6426
rect 515904 -7654 516504 -6662
rect 533904 -7066 534504 31158
rect 540804 704838 541404 705830
rect 540804 704602 540986 704838
rect 541222 704602 541404 704838
rect 540804 704518 541404 704602
rect 540804 704282 540986 704518
rect 541222 704282 541404 704518
rect 540804 686294 541404 704282
rect 540804 686058 540986 686294
rect 541222 686058 541404 686294
rect 540804 650294 541404 686058
rect 540804 650058 540986 650294
rect 541222 650058 541404 650294
rect 540804 614294 541404 650058
rect 540804 614058 540986 614294
rect 541222 614058 541404 614294
rect 540804 578294 541404 614058
rect 540804 578058 540986 578294
rect 541222 578058 541404 578294
rect 540804 542294 541404 578058
rect 540804 542058 540986 542294
rect 541222 542058 541404 542294
rect 540804 506294 541404 542058
rect 540804 506058 540986 506294
rect 541222 506058 541404 506294
rect 540804 470294 541404 506058
rect 540804 470058 540986 470294
rect 541222 470058 541404 470294
rect 540804 434294 541404 470058
rect 540804 434058 540986 434294
rect 541222 434058 541404 434294
rect 540804 398294 541404 434058
rect 540804 398058 540986 398294
rect 541222 398058 541404 398294
rect 540804 362294 541404 398058
rect 540804 362058 540986 362294
rect 541222 362058 541404 362294
rect 540804 326294 541404 362058
rect 540804 326058 540986 326294
rect 541222 326058 541404 326294
rect 540804 290294 541404 326058
rect 540804 290058 540986 290294
rect 541222 290058 541404 290294
rect 540804 254294 541404 290058
rect 540804 254058 540986 254294
rect 541222 254058 541404 254294
rect 540804 218294 541404 254058
rect 540804 218058 540986 218294
rect 541222 218058 541404 218294
rect 540804 182294 541404 218058
rect 540804 182058 540986 182294
rect 541222 182058 541404 182294
rect 540804 146294 541404 182058
rect 540804 146058 540986 146294
rect 541222 146058 541404 146294
rect 540804 110294 541404 146058
rect 540804 110058 540986 110294
rect 541222 110058 541404 110294
rect 540804 74294 541404 110058
rect 540804 74058 540986 74294
rect 541222 74058 541404 74294
rect 540804 38294 541404 74058
rect 540804 38058 540986 38294
rect 541222 38058 541404 38294
rect 540804 2294 541404 38058
rect 540804 2058 540986 2294
rect 541222 2058 541404 2294
rect 540804 -346 541404 2058
rect 540804 -582 540986 -346
rect 541222 -582 541404 -346
rect 540804 -666 541404 -582
rect 540804 -902 540986 -666
rect 541222 -902 541404 -666
rect 540804 -1894 541404 -902
rect 544504 689994 545104 706202
rect 544504 689758 544686 689994
rect 544922 689758 545104 689994
rect 544504 653994 545104 689758
rect 544504 653758 544686 653994
rect 544922 653758 545104 653994
rect 544504 617994 545104 653758
rect 544504 617758 544686 617994
rect 544922 617758 545104 617994
rect 544504 581994 545104 617758
rect 544504 581758 544686 581994
rect 544922 581758 545104 581994
rect 544504 545994 545104 581758
rect 544504 545758 544686 545994
rect 544922 545758 545104 545994
rect 544504 509994 545104 545758
rect 544504 509758 544686 509994
rect 544922 509758 545104 509994
rect 544504 473994 545104 509758
rect 544504 473758 544686 473994
rect 544922 473758 545104 473994
rect 544504 437994 545104 473758
rect 544504 437758 544686 437994
rect 544922 437758 545104 437994
rect 544504 401994 545104 437758
rect 544504 401758 544686 401994
rect 544922 401758 545104 401994
rect 544504 365994 545104 401758
rect 544504 365758 544686 365994
rect 544922 365758 545104 365994
rect 544504 329994 545104 365758
rect 544504 329758 544686 329994
rect 544922 329758 545104 329994
rect 544504 293994 545104 329758
rect 544504 293758 544686 293994
rect 544922 293758 545104 293994
rect 544504 257994 545104 293758
rect 544504 257758 544686 257994
rect 544922 257758 545104 257994
rect 544504 221994 545104 257758
rect 544504 221758 544686 221994
rect 544922 221758 545104 221994
rect 544504 185994 545104 221758
rect 544504 185758 544686 185994
rect 544922 185758 545104 185994
rect 544504 149994 545104 185758
rect 544504 149758 544686 149994
rect 544922 149758 545104 149994
rect 544504 113994 545104 149758
rect 544504 113758 544686 113994
rect 544922 113758 545104 113994
rect 544504 77994 545104 113758
rect 544504 77758 544686 77994
rect 544922 77758 545104 77994
rect 544504 41994 545104 77758
rect 544504 41758 544686 41994
rect 544922 41758 545104 41994
rect 544504 5994 545104 41758
rect 544504 5758 544686 5994
rect 544922 5758 545104 5994
rect 544504 -2266 545104 5758
rect 544504 -2502 544686 -2266
rect 544922 -2502 545104 -2266
rect 544504 -2586 545104 -2502
rect 544504 -2822 544686 -2586
rect 544922 -2822 545104 -2586
rect 544504 -3814 545104 -2822
rect 548204 693694 548804 708122
rect 548204 693458 548386 693694
rect 548622 693458 548804 693694
rect 548204 657694 548804 693458
rect 548204 657458 548386 657694
rect 548622 657458 548804 657694
rect 548204 621694 548804 657458
rect 548204 621458 548386 621694
rect 548622 621458 548804 621694
rect 548204 585694 548804 621458
rect 548204 585458 548386 585694
rect 548622 585458 548804 585694
rect 548204 549694 548804 585458
rect 548204 549458 548386 549694
rect 548622 549458 548804 549694
rect 548204 513694 548804 549458
rect 548204 513458 548386 513694
rect 548622 513458 548804 513694
rect 548204 477694 548804 513458
rect 548204 477458 548386 477694
rect 548622 477458 548804 477694
rect 548204 441694 548804 477458
rect 548204 441458 548386 441694
rect 548622 441458 548804 441694
rect 548204 405694 548804 441458
rect 548204 405458 548386 405694
rect 548622 405458 548804 405694
rect 548204 369694 548804 405458
rect 548204 369458 548386 369694
rect 548622 369458 548804 369694
rect 548204 333694 548804 369458
rect 548204 333458 548386 333694
rect 548622 333458 548804 333694
rect 548204 297694 548804 333458
rect 548204 297458 548386 297694
rect 548622 297458 548804 297694
rect 548204 261694 548804 297458
rect 548204 261458 548386 261694
rect 548622 261458 548804 261694
rect 548204 225694 548804 261458
rect 548204 225458 548386 225694
rect 548622 225458 548804 225694
rect 548204 189694 548804 225458
rect 548204 189458 548386 189694
rect 548622 189458 548804 189694
rect 548204 153694 548804 189458
rect 548204 153458 548386 153694
rect 548622 153458 548804 153694
rect 548204 117694 548804 153458
rect 548204 117458 548386 117694
rect 548622 117458 548804 117694
rect 548204 81694 548804 117458
rect 548204 81458 548386 81694
rect 548622 81458 548804 81694
rect 548204 45694 548804 81458
rect 548204 45458 548386 45694
rect 548622 45458 548804 45694
rect 548204 9694 548804 45458
rect 548204 9458 548386 9694
rect 548622 9458 548804 9694
rect 548204 -4186 548804 9458
rect 548204 -4422 548386 -4186
rect 548622 -4422 548804 -4186
rect 548204 -4506 548804 -4422
rect 548204 -4742 548386 -4506
rect 548622 -4742 548804 -4506
rect 548204 -5734 548804 -4742
rect 551904 697394 552504 710042
rect 569904 711558 570504 711590
rect 569904 711322 570086 711558
rect 570322 711322 570504 711558
rect 569904 711238 570504 711322
rect 569904 711002 570086 711238
rect 570322 711002 570504 711238
rect 566204 709638 566804 709670
rect 566204 709402 566386 709638
rect 566622 709402 566804 709638
rect 566204 709318 566804 709402
rect 566204 709082 566386 709318
rect 566622 709082 566804 709318
rect 562504 707718 563104 707750
rect 562504 707482 562686 707718
rect 562922 707482 563104 707718
rect 562504 707398 563104 707482
rect 562504 707162 562686 707398
rect 562922 707162 563104 707398
rect 551904 697158 552086 697394
rect 552322 697158 552504 697394
rect 551904 661394 552504 697158
rect 551904 661158 552086 661394
rect 552322 661158 552504 661394
rect 551904 625394 552504 661158
rect 551904 625158 552086 625394
rect 552322 625158 552504 625394
rect 551904 589394 552504 625158
rect 551904 589158 552086 589394
rect 552322 589158 552504 589394
rect 551904 553394 552504 589158
rect 551904 553158 552086 553394
rect 552322 553158 552504 553394
rect 551904 517394 552504 553158
rect 551904 517158 552086 517394
rect 552322 517158 552504 517394
rect 551904 481394 552504 517158
rect 551904 481158 552086 481394
rect 552322 481158 552504 481394
rect 551904 445394 552504 481158
rect 551904 445158 552086 445394
rect 552322 445158 552504 445394
rect 551904 409394 552504 445158
rect 551904 409158 552086 409394
rect 552322 409158 552504 409394
rect 551904 373394 552504 409158
rect 551904 373158 552086 373394
rect 552322 373158 552504 373394
rect 551904 337394 552504 373158
rect 551904 337158 552086 337394
rect 552322 337158 552504 337394
rect 551904 301394 552504 337158
rect 551904 301158 552086 301394
rect 552322 301158 552504 301394
rect 551904 265394 552504 301158
rect 551904 265158 552086 265394
rect 552322 265158 552504 265394
rect 551904 229394 552504 265158
rect 551904 229158 552086 229394
rect 552322 229158 552504 229394
rect 551904 193394 552504 229158
rect 551904 193158 552086 193394
rect 552322 193158 552504 193394
rect 551904 157394 552504 193158
rect 551904 157158 552086 157394
rect 552322 157158 552504 157394
rect 551904 121394 552504 157158
rect 551904 121158 552086 121394
rect 552322 121158 552504 121394
rect 551904 85394 552504 121158
rect 551904 85158 552086 85394
rect 552322 85158 552504 85394
rect 551904 49394 552504 85158
rect 551904 49158 552086 49394
rect 552322 49158 552504 49394
rect 551904 13394 552504 49158
rect 551904 13158 552086 13394
rect 552322 13158 552504 13394
rect 533904 -7302 534086 -7066
rect 534322 -7302 534504 -7066
rect 533904 -7386 534504 -7302
rect 533904 -7622 534086 -7386
rect 534322 -7622 534504 -7386
rect 533904 -7654 534504 -7622
rect 551904 -6106 552504 13158
rect 558804 705798 559404 705830
rect 558804 705562 558986 705798
rect 559222 705562 559404 705798
rect 558804 705478 559404 705562
rect 558804 705242 558986 705478
rect 559222 705242 559404 705478
rect 558804 668294 559404 705242
rect 558804 668058 558986 668294
rect 559222 668058 559404 668294
rect 558804 632294 559404 668058
rect 558804 632058 558986 632294
rect 559222 632058 559404 632294
rect 558804 596294 559404 632058
rect 558804 596058 558986 596294
rect 559222 596058 559404 596294
rect 558804 560294 559404 596058
rect 558804 560058 558986 560294
rect 559222 560058 559404 560294
rect 558804 524294 559404 560058
rect 558804 524058 558986 524294
rect 559222 524058 559404 524294
rect 558804 488294 559404 524058
rect 558804 488058 558986 488294
rect 559222 488058 559404 488294
rect 558804 452294 559404 488058
rect 558804 452058 558986 452294
rect 559222 452058 559404 452294
rect 558804 416294 559404 452058
rect 558804 416058 558986 416294
rect 559222 416058 559404 416294
rect 558804 380294 559404 416058
rect 558804 380058 558986 380294
rect 559222 380058 559404 380294
rect 558804 344294 559404 380058
rect 558804 344058 558986 344294
rect 559222 344058 559404 344294
rect 558804 308294 559404 344058
rect 558804 308058 558986 308294
rect 559222 308058 559404 308294
rect 558804 272294 559404 308058
rect 558804 272058 558986 272294
rect 559222 272058 559404 272294
rect 558804 236294 559404 272058
rect 558804 236058 558986 236294
rect 559222 236058 559404 236294
rect 558804 200294 559404 236058
rect 558804 200058 558986 200294
rect 559222 200058 559404 200294
rect 558804 164294 559404 200058
rect 558804 164058 558986 164294
rect 559222 164058 559404 164294
rect 558804 128294 559404 164058
rect 558804 128058 558986 128294
rect 559222 128058 559404 128294
rect 558804 92294 559404 128058
rect 558804 92058 558986 92294
rect 559222 92058 559404 92294
rect 558804 56294 559404 92058
rect 558804 56058 558986 56294
rect 559222 56058 559404 56294
rect 558804 20294 559404 56058
rect 558804 20058 558986 20294
rect 559222 20058 559404 20294
rect 558804 -1306 559404 20058
rect 558804 -1542 558986 -1306
rect 559222 -1542 559404 -1306
rect 558804 -1626 559404 -1542
rect 558804 -1862 558986 -1626
rect 559222 -1862 559404 -1626
rect 558804 -1894 559404 -1862
rect 562504 671994 563104 707162
rect 562504 671758 562686 671994
rect 562922 671758 563104 671994
rect 562504 635994 563104 671758
rect 562504 635758 562686 635994
rect 562922 635758 563104 635994
rect 562504 599994 563104 635758
rect 562504 599758 562686 599994
rect 562922 599758 563104 599994
rect 562504 563994 563104 599758
rect 562504 563758 562686 563994
rect 562922 563758 563104 563994
rect 562504 527994 563104 563758
rect 562504 527758 562686 527994
rect 562922 527758 563104 527994
rect 562504 491994 563104 527758
rect 562504 491758 562686 491994
rect 562922 491758 563104 491994
rect 562504 455994 563104 491758
rect 562504 455758 562686 455994
rect 562922 455758 563104 455994
rect 562504 419994 563104 455758
rect 562504 419758 562686 419994
rect 562922 419758 563104 419994
rect 562504 383994 563104 419758
rect 562504 383758 562686 383994
rect 562922 383758 563104 383994
rect 562504 347994 563104 383758
rect 562504 347758 562686 347994
rect 562922 347758 563104 347994
rect 562504 311994 563104 347758
rect 562504 311758 562686 311994
rect 562922 311758 563104 311994
rect 562504 275994 563104 311758
rect 562504 275758 562686 275994
rect 562922 275758 563104 275994
rect 562504 239994 563104 275758
rect 562504 239758 562686 239994
rect 562922 239758 563104 239994
rect 562504 203994 563104 239758
rect 562504 203758 562686 203994
rect 562922 203758 563104 203994
rect 562504 167994 563104 203758
rect 562504 167758 562686 167994
rect 562922 167758 563104 167994
rect 562504 131994 563104 167758
rect 562504 131758 562686 131994
rect 562922 131758 563104 131994
rect 562504 95994 563104 131758
rect 562504 95758 562686 95994
rect 562922 95758 563104 95994
rect 562504 59994 563104 95758
rect 562504 59758 562686 59994
rect 562922 59758 563104 59994
rect 562504 23994 563104 59758
rect 562504 23758 562686 23994
rect 562922 23758 563104 23994
rect 562504 -3226 563104 23758
rect 562504 -3462 562686 -3226
rect 562922 -3462 563104 -3226
rect 562504 -3546 563104 -3462
rect 562504 -3782 562686 -3546
rect 562922 -3782 563104 -3546
rect 562504 -3814 563104 -3782
rect 566204 675694 566804 709082
rect 566204 675458 566386 675694
rect 566622 675458 566804 675694
rect 566204 639694 566804 675458
rect 566204 639458 566386 639694
rect 566622 639458 566804 639694
rect 566204 603694 566804 639458
rect 566204 603458 566386 603694
rect 566622 603458 566804 603694
rect 566204 567694 566804 603458
rect 566204 567458 566386 567694
rect 566622 567458 566804 567694
rect 566204 531694 566804 567458
rect 566204 531458 566386 531694
rect 566622 531458 566804 531694
rect 566204 495694 566804 531458
rect 566204 495458 566386 495694
rect 566622 495458 566804 495694
rect 566204 459694 566804 495458
rect 566204 459458 566386 459694
rect 566622 459458 566804 459694
rect 566204 423694 566804 459458
rect 566204 423458 566386 423694
rect 566622 423458 566804 423694
rect 566204 387694 566804 423458
rect 566204 387458 566386 387694
rect 566622 387458 566804 387694
rect 566204 351694 566804 387458
rect 566204 351458 566386 351694
rect 566622 351458 566804 351694
rect 566204 315694 566804 351458
rect 566204 315458 566386 315694
rect 566622 315458 566804 315694
rect 566204 279694 566804 315458
rect 566204 279458 566386 279694
rect 566622 279458 566804 279694
rect 566204 243694 566804 279458
rect 566204 243458 566386 243694
rect 566622 243458 566804 243694
rect 566204 207694 566804 243458
rect 566204 207458 566386 207694
rect 566622 207458 566804 207694
rect 566204 171694 566804 207458
rect 566204 171458 566386 171694
rect 566622 171458 566804 171694
rect 566204 135694 566804 171458
rect 566204 135458 566386 135694
rect 566622 135458 566804 135694
rect 566204 99694 566804 135458
rect 566204 99458 566386 99694
rect 566622 99458 566804 99694
rect 566204 63694 566804 99458
rect 566204 63458 566386 63694
rect 566622 63458 566804 63694
rect 566204 27694 566804 63458
rect 566204 27458 566386 27694
rect 566622 27458 566804 27694
rect 566204 -5146 566804 27458
rect 566204 -5382 566386 -5146
rect 566622 -5382 566804 -5146
rect 566204 -5466 566804 -5382
rect 566204 -5702 566386 -5466
rect 566622 -5702 566804 -5466
rect 566204 -5734 566804 -5702
rect 569904 679394 570504 711002
rect 592030 711558 592650 711590
rect 592030 711322 592062 711558
rect 592298 711322 592382 711558
rect 592618 711322 592650 711558
rect 592030 711238 592650 711322
rect 592030 711002 592062 711238
rect 592298 711002 592382 711238
rect 592618 711002 592650 711238
rect 591070 710598 591690 710630
rect 591070 710362 591102 710598
rect 591338 710362 591422 710598
rect 591658 710362 591690 710598
rect 591070 710278 591690 710362
rect 591070 710042 591102 710278
rect 591338 710042 591422 710278
rect 591658 710042 591690 710278
rect 590110 709638 590730 709670
rect 590110 709402 590142 709638
rect 590378 709402 590462 709638
rect 590698 709402 590730 709638
rect 590110 709318 590730 709402
rect 590110 709082 590142 709318
rect 590378 709082 590462 709318
rect 590698 709082 590730 709318
rect 589150 708678 589770 708710
rect 589150 708442 589182 708678
rect 589418 708442 589502 708678
rect 589738 708442 589770 708678
rect 589150 708358 589770 708442
rect 589150 708122 589182 708358
rect 589418 708122 589502 708358
rect 589738 708122 589770 708358
rect 580504 706758 581104 707750
rect 588190 707718 588810 707750
rect 588190 707482 588222 707718
rect 588458 707482 588542 707718
rect 588778 707482 588810 707718
rect 588190 707398 588810 707482
rect 588190 707162 588222 707398
rect 588458 707162 588542 707398
rect 588778 707162 588810 707398
rect 580504 706522 580686 706758
rect 580922 706522 581104 706758
rect 580504 706438 581104 706522
rect 580504 706202 580686 706438
rect 580922 706202 581104 706438
rect 569904 679158 570086 679394
rect 570322 679158 570504 679394
rect 569904 643394 570504 679158
rect 569904 643158 570086 643394
rect 570322 643158 570504 643394
rect 569904 607394 570504 643158
rect 569904 607158 570086 607394
rect 570322 607158 570504 607394
rect 569904 571394 570504 607158
rect 569904 571158 570086 571394
rect 570322 571158 570504 571394
rect 569904 535394 570504 571158
rect 569904 535158 570086 535394
rect 570322 535158 570504 535394
rect 569904 499394 570504 535158
rect 569904 499158 570086 499394
rect 570322 499158 570504 499394
rect 569904 463394 570504 499158
rect 569904 463158 570086 463394
rect 570322 463158 570504 463394
rect 569904 427394 570504 463158
rect 569904 427158 570086 427394
rect 570322 427158 570504 427394
rect 569904 391394 570504 427158
rect 569904 391158 570086 391394
rect 570322 391158 570504 391394
rect 569904 355394 570504 391158
rect 569904 355158 570086 355394
rect 570322 355158 570504 355394
rect 569904 319394 570504 355158
rect 569904 319158 570086 319394
rect 570322 319158 570504 319394
rect 569904 283394 570504 319158
rect 569904 283158 570086 283394
rect 570322 283158 570504 283394
rect 569904 247394 570504 283158
rect 569904 247158 570086 247394
rect 570322 247158 570504 247394
rect 569904 211394 570504 247158
rect 569904 211158 570086 211394
rect 570322 211158 570504 211394
rect 569904 175394 570504 211158
rect 569904 175158 570086 175394
rect 570322 175158 570504 175394
rect 569904 139394 570504 175158
rect 569904 139158 570086 139394
rect 570322 139158 570504 139394
rect 569904 103394 570504 139158
rect 569904 103158 570086 103394
rect 570322 103158 570504 103394
rect 569904 67394 570504 103158
rect 569904 67158 570086 67394
rect 570322 67158 570504 67394
rect 569904 31394 570504 67158
rect 569904 31158 570086 31394
rect 570322 31158 570504 31394
rect 551904 -6342 552086 -6106
rect 552322 -6342 552504 -6106
rect 551904 -6426 552504 -6342
rect 551904 -6662 552086 -6426
rect 552322 -6662 552504 -6426
rect 551904 -7654 552504 -6662
rect 569904 -7066 570504 31158
rect 576804 704838 577404 705830
rect 576804 704602 576986 704838
rect 577222 704602 577404 704838
rect 576804 704518 577404 704602
rect 576804 704282 576986 704518
rect 577222 704282 577404 704518
rect 576804 686294 577404 704282
rect 576804 686058 576986 686294
rect 577222 686058 577404 686294
rect 576804 650294 577404 686058
rect 576804 650058 576986 650294
rect 577222 650058 577404 650294
rect 576804 614294 577404 650058
rect 576804 614058 576986 614294
rect 577222 614058 577404 614294
rect 576804 578294 577404 614058
rect 576804 578058 576986 578294
rect 577222 578058 577404 578294
rect 576804 542294 577404 578058
rect 576804 542058 576986 542294
rect 577222 542058 577404 542294
rect 576804 506294 577404 542058
rect 576804 506058 576986 506294
rect 577222 506058 577404 506294
rect 576804 470294 577404 506058
rect 576804 470058 576986 470294
rect 577222 470058 577404 470294
rect 576804 434294 577404 470058
rect 576804 434058 576986 434294
rect 577222 434058 577404 434294
rect 576804 398294 577404 434058
rect 576804 398058 576986 398294
rect 577222 398058 577404 398294
rect 576804 362294 577404 398058
rect 576804 362058 576986 362294
rect 577222 362058 577404 362294
rect 576804 326294 577404 362058
rect 576804 326058 576986 326294
rect 577222 326058 577404 326294
rect 576804 290294 577404 326058
rect 576804 290058 576986 290294
rect 577222 290058 577404 290294
rect 576804 254294 577404 290058
rect 576804 254058 576986 254294
rect 577222 254058 577404 254294
rect 576804 218294 577404 254058
rect 576804 218058 576986 218294
rect 577222 218058 577404 218294
rect 576804 182294 577404 218058
rect 576804 182058 576986 182294
rect 577222 182058 577404 182294
rect 576804 146294 577404 182058
rect 576804 146058 576986 146294
rect 577222 146058 577404 146294
rect 576804 110294 577404 146058
rect 576804 110058 576986 110294
rect 577222 110058 577404 110294
rect 576804 74294 577404 110058
rect 576804 74058 576986 74294
rect 577222 74058 577404 74294
rect 576804 38294 577404 74058
rect 576804 38058 576986 38294
rect 577222 38058 577404 38294
rect 576804 2294 577404 38058
rect 576804 2058 576986 2294
rect 577222 2058 577404 2294
rect 576804 -346 577404 2058
rect 576804 -582 576986 -346
rect 577222 -582 577404 -346
rect 576804 -666 577404 -582
rect 576804 -902 576986 -666
rect 577222 -902 577404 -666
rect 576804 -1894 577404 -902
rect 580504 689994 581104 706202
rect 587230 706758 587850 706790
rect 587230 706522 587262 706758
rect 587498 706522 587582 706758
rect 587818 706522 587850 706758
rect 587230 706438 587850 706522
rect 587230 706202 587262 706438
rect 587498 706202 587582 706438
rect 587818 706202 587850 706438
rect 586270 705798 586890 705830
rect 586270 705562 586302 705798
rect 586538 705562 586622 705798
rect 586858 705562 586890 705798
rect 586270 705478 586890 705562
rect 586270 705242 586302 705478
rect 586538 705242 586622 705478
rect 586858 705242 586890 705478
rect 580504 689758 580686 689994
rect 580922 689758 581104 689994
rect 580504 653994 581104 689758
rect 580504 653758 580686 653994
rect 580922 653758 581104 653994
rect 580504 617994 581104 653758
rect 580504 617758 580686 617994
rect 580922 617758 581104 617994
rect 580504 581994 581104 617758
rect 580504 581758 580686 581994
rect 580922 581758 581104 581994
rect 580504 545994 581104 581758
rect 580504 545758 580686 545994
rect 580922 545758 581104 545994
rect 580504 509994 581104 545758
rect 580504 509758 580686 509994
rect 580922 509758 581104 509994
rect 580504 473994 581104 509758
rect 580504 473758 580686 473994
rect 580922 473758 581104 473994
rect 580504 437994 581104 473758
rect 580504 437758 580686 437994
rect 580922 437758 581104 437994
rect 580504 401994 581104 437758
rect 580504 401758 580686 401994
rect 580922 401758 581104 401994
rect 580504 365994 581104 401758
rect 580504 365758 580686 365994
rect 580922 365758 581104 365994
rect 580504 329994 581104 365758
rect 580504 329758 580686 329994
rect 580922 329758 581104 329994
rect 580504 293994 581104 329758
rect 580504 293758 580686 293994
rect 580922 293758 581104 293994
rect 580504 257994 581104 293758
rect 580504 257758 580686 257994
rect 580922 257758 581104 257994
rect 580504 221994 581104 257758
rect 580504 221758 580686 221994
rect 580922 221758 581104 221994
rect 580504 185994 581104 221758
rect 580504 185758 580686 185994
rect 580922 185758 581104 185994
rect 580504 149994 581104 185758
rect 580504 149758 580686 149994
rect 580922 149758 581104 149994
rect 580504 113994 581104 149758
rect 580504 113758 580686 113994
rect 580922 113758 581104 113994
rect 580504 77994 581104 113758
rect 580504 77758 580686 77994
rect 580922 77758 581104 77994
rect 580504 41994 581104 77758
rect 580504 41758 580686 41994
rect 580922 41758 581104 41994
rect 580504 5994 581104 41758
rect 580504 5758 580686 5994
rect 580922 5758 581104 5994
rect 580504 -2266 581104 5758
rect 585310 704838 585930 704870
rect 585310 704602 585342 704838
rect 585578 704602 585662 704838
rect 585898 704602 585930 704838
rect 585310 704518 585930 704602
rect 585310 704282 585342 704518
rect 585578 704282 585662 704518
rect 585898 704282 585930 704518
rect 585310 686294 585930 704282
rect 585310 686058 585342 686294
rect 585578 686058 585662 686294
rect 585898 686058 585930 686294
rect 585310 650294 585930 686058
rect 585310 650058 585342 650294
rect 585578 650058 585662 650294
rect 585898 650058 585930 650294
rect 585310 614294 585930 650058
rect 585310 614058 585342 614294
rect 585578 614058 585662 614294
rect 585898 614058 585930 614294
rect 585310 578294 585930 614058
rect 585310 578058 585342 578294
rect 585578 578058 585662 578294
rect 585898 578058 585930 578294
rect 585310 542294 585930 578058
rect 585310 542058 585342 542294
rect 585578 542058 585662 542294
rect 585898 542058 585930 542294
rect 585310 506294 585930 542058
rect 585310 506058 585342 506294
rect 585578 506058 585662 506294
rect 585898 506058 585930 506294
rect 585310 470294 585930 506058
rect 585310 470058 585342 470294
rect 585578 470058 585662 470294
rect 585898 470058 585930 470294
rect 585310 434294 585930 470058
rect 585310 434058 585342 434294
rect 585578 434058 585662 434294
rect 585898 434058 585930 434294
rect 585310 398294 585930 434058
rect 585310 398058 585342 398294
rect 585578 398058 585662 398294
rect 585898 398058 585930 398294
rect 585310 362294 585930 398058
rect 585310 362058 585342 362294
rect 585578 362058 585662 362294
rect 585898 362058 585930 362294
rect 585310 326294 585930 362058
rect 585310 326058 585342 326294
rect 585578 326058 585662 326294
rect 585898 326058 585930 326294
rect 585310 290294 585930 326058
rect 585310 290058 585342 290294
rect 585578 290058 585662 290294
rect 585898 290058 585930 290294
rect 585310 254294 585930 290058
rect 585310 254058 585342 254294
rect 585578 254058 585662 254294
rect 585898 254058 585930 254294
rect 585310 218294 585930 254058
rect 585310 218058 585342 218294
rect 585578 218058 585662 218294
rect 585898 218058 585930 218294
rect 585310 182294 585930 218058
rect 585310 182058 585342 182294
rect 585578 182058 585662 182294
rect 585898 182058 585930 182294
rect 585310 146294 585930 182058
rect 585310 146058 585342 146294
rect 585578 146058 585662 146294
rect 585898 146058 585930 146294
rect 585310 110294 585930 146058
rect 585310 110058 585342 110294
rect 585578 110058 585662 110294
rect 585898 110058 585930 110294
rect 585310 74294 585930 110058
rect 585310 74058 585342 74294
rect 585578 74058 585662 74294
rect 585898 74058 585930 74294
rect 585310 38294 585930 74058
rect 585310 38058 585342 38294
rect 585578 38058 585662 38294
rect 585898 38058 585930 38294
rect 585310 2294 585930 38058
rect 585310 2058 585342 2294
rect 585578 2058 585662 2294
rect 585898 2058 585930 2294
rect 585310 -346 585930 2058
rect 585310 -582 585342 -346
rect 585578 -582 585662 -346
rect 585898 -582 585930 -346
rect 585310 -666 585930 -582
rect 585310 -902 585342 -666
rect 585578 -902 585662 -666
rect 585898 -902 585930 -666
rect 585310 -934 585930 -902
rect 586270 668294 586890 705242
rect 586270 668058 586302 668294
rect 586538 668058 586622 668294
rect 586858 668058 586890 668294
rect 586270 632294 586890 668058
rect 586270 632058 586302 632294
rect 586538 632058 586622 632294
rect 586858 632058 586890 632294
rect 586270 596294 586890 632058
rect 586270 596058 586302 596294
rect 586538 596058 586622 596294
rect 586858 596058 586890 596294
rect 586270 560294 586890 596058
rect 586270 560058 586302 560294
rect 586538 560058 586622 560294
rect 586858 560058 586890 560294
rect 586270 524294 586890 560058
rect 586270 524058 586302 524294
rect 586538 524058 586622 524294
rect 586858 524058 586890 524294
rect 586270 488294 586890 524058
rect 586270 488058 586302 488294
rect 586538 488058 586622 488294
rect 586858 488058 586890 488294
rect 586270 452294 586890 488058
rect 586270 452058 586302 452294
rect 586538 452058 586622 452294
rect 586858 452058 586890 452294
rect 586270 416294 586890 452058
rect 586270 416058 586302 416294
rect 586538 416058 586622 416294
rect 586858 416058 586890 416294
rect 586270 380294 586890 416058
rect 586270 380058 586302 380294
rect 586538 380058 586622 380294
rect 586858 380058 586890 380294
rect 586270 344294 586890 380058
rect 586270 344058 586302 344294
rect 586538 344058 586622 344294
rect 586858 344058 586890 344294
rect 586270 308294 586890 344058
rect 586270 308058 586302 308294
rect 586538 308058 586622 308294
rect 586858 308058 586890 308294
rect 586270 272294 586890 308058
rect 586270 272058 586302 272294
rect 586538 272058 586622 272294
rect 586858 272058 586890 272294
rect 586270 236294 586890 272058
rect 586270 236058 586302 236294
rect 586538 236058 586622 236294
rect 586858 236058 586890 236294
rect 586270 200294 586890 236058
rect 586270 200058 586302 200294
rect 586538 200058 586622 200294
rect 586858 200058 586890 200294
rect 586270 164294 586890 200058
rect 586270 164058 586302 164294
rect 586538 164058 586622 164294
rect 586858 164058 586890 164294
rect 586270 128294 586890 164058
rect 586270 128058 586302 128294
rect 586538 128058 586622 128294
rect 586858 128058 586890 128294
rect 586270 92294 586890 128058
rect 586270 92058 586302 92294
rect 586538 92058 586622 92294
rect 586858 92058 586890 92294
rect 586270 56294 586890 92058
rect 586270 56058 586302 56294
rect 586538 56058 586622 56294
rect 586858 56058 586890 56294
rect 586270 20294 586890 56058
rect 586270 20058 586302 20294
rect 586538 20058 586622 20294
rect 586858 20058 586890 20294
rect 586270 -1306 586890 20058
rect 586270 -1542 586302 -1306
rect 586538 -1542 586622 -1306
rect 586858 -1542 586890 -1306
rect 586270 -1626 586890 -1542
rect 586270 -1862 586302 -1626
rect 586538 -1862 586622 -1626
rect 586858 -1862 586890 -1626
rect 586270 -1894 586890 -1862
rect 587230 689994 587850 706202
rect 587230 689758 587262 689994
rect 587498 689758 587582 689994
rect 587818 689758 587850 689994
rect 587230 653994 587850 689758
rect 587230 653758 587262 653994
rect 587498 653758 587582 653994
rect 587818 653758 587850 653994
rect 587230 617994 587850 653758
rect 587230 617758 587262 617994
rect 587498 617758 587582 617994
rect 587818 617758 587850 617994
rect 587230 581994 587850 617758
rect 587230 581758 587262 581994
rect 587498 581758 587582 581994
rect 587818 581758 587850 581994
rect 587230 545994 587850 581758
rect 587230 545758 587262 545994
rect 587498 545758 587582 545994
rect 587818 545758 587850 545994
rect 587230 509994 587850 545758
rect 587230 509758 587262 509994
rect 587498 509758 587582 509994
rect 587818 509758 587850 509994
rect 587230 473994 587850 509758
rect 587230 473758 587262 473994
rect 587498 473758 587582 473994
rect 587818 473758 587850 473994
rect 587230 437994 587850 473758
rect 587230 437758 587262 437994
rect 587498 437758 587582 437994
rect 587818 437758 587850 437994
rect 587230 401994 587850 437758
rect 587230 401758 587262 401994
rect 587498 401758 587582 401994
rect 587818 401758 587850 401994
rect 587230 365994 587850 401758
rect 587230 365758 587262 365994
rect 587498 365758 587582 365994
rect 587818 365758 587850 365994
rect 587230 329994 587850 365758
rect 587230 329758 587262 329994
rect 587498 329758 587582 329994
rect 587818 329758 587850 329994
rect 587230 293994 587850 329758
rect 587230 293758 587262 293994
rect 587498 293758 587582 293994
rect 587818 293758 587850 293994
rect 587230 257994 587850 293758
rect 587230 257758 587262 257994
rect 587498 257758 587582 257994
rect 587818 257758 587850 257994
rect 587230 221994 587850 257758
rect 587230 221758 587262 221994
rect 587498 221758 587582 221994
rect 587818 221758 587850 221994
rect 587230 185994 587850 221758
rect 587230 185758 587262 185994
rect 587498 185758 587582 185994
rect 587818 185758 587850 185994
rect 587230 149994 587850 185758
rect 587230 149758 587262 149994
rect 587498 149758 587582 149994
rect 587818 149758 587850 149994
rect 587230 113994 587850 149758
rect 587230 113758 587262 113994
rect 587498 113758 587582 113994
rect 587818 113758 587850 113994
rect 587230 77994 587850 113758
rect 587230 77758 587262 77994
rect 587498 77758 587582 77994
rect 587818 77758 587850 77994
rect 587230 41994 587850 77758
rect 587230 41758 587262 41994
rect 587498 41758 587582 41994
rect 587818 41758 587850 41994
rect 587230 5994 587850 41758
rect 587230 5758 587262 5994
rect 587498 5758 587582 5994
rect 587818 5758 587850 5994
rect 580504 -2502 580686 -2266
rect 580922 -2502 581104 -2266
rect 580504 -2586 581104 -2502
rect 580504 -2822 580686 -2586
rect 580922 -2822 581104 -2586
rect 580504 -3814 581104 -2822
rect 587230 -2266 587850 5758
rect 587230 -2502 587262 -2266
rect 587498 -2502 587582 -2266
rect 587818 -2502 587850 -2266
rect 587230 -2586 587850 -2502
rect 587230 -2822 587262 -2586
rect 587498 -2822 587582 -2586
rect 587818 -2822 587850 -2586
rect 587230 -2854 587850 -2822
rect 588190 671994 588810 707162
rect 588190 671758 588222 671994
rect 588458 671758 588542 671994
rect 588778 671758 588810 671994
rect 588190 635994 588810 671758
rect 588190 635758 588222 635994
rect 588458 635758 588542 635994
rect 588778 635758 588810 635994
rect 588190 599994 588810 635758
rect 588190 599758 588222 599994
rect 588458 599758 588542 599994
rect 588778 599758 588810 599994
rect 588190 563994 588810 599758
rect 588190 563758 588222 563994
rect 588458 563758 588542 563994
rect 588778 563758 588810 563994
rect 588190 527994 588810 563758
rect 588190 527758 588222 527994
rect 588458 527758 588542 527994
rect 588778 527758 588810 527994
rect 588190 491994 588810 527758
rect 588190 491758 588222 491994
rect 588458 491758 588542 491994
rect 588778 491758 588810 491994
rect 588190 455994 588810 491758
rect 588190 455758 588222 455994
rect 588458 455758 588542 455994
rect 588778 455758 588810 455994
rect 588190 419994 588810 455758
rect 588190 419758 588222 419994
rect 588458 419758 588542 419994
rect 588778 419758 588810 419994
rect 588190 383994 588810 419758
rect 588190 383758 588222 383994
rect 588458 383758 588542 383994
rect 588778 383758 588810 383994
rect 588190 347994 588810 383758
rect 588190 347758 588222 347994
rect 588458 347758 588542 347994
rect 588778 347758 588810 347994
rect 588190 311994 588810 347758
rect 588190 311758 588222 311994
rect 588458 311758 588542 311994
rect 588778 311758 588810 311994
rect 588190 275994 588810 311758
rect 588190 275758 588222 275994
rect 588458 275758 588542 275994
rect 588778 275758 588810 275994
rect 588190 239994 588810 275758
rect 588190 239758 588222 239994
rect 588458 239758 588542 239994
rect 588778 239758 588810 239994
rect 588190 203994 588810 239758
rect 588190 203758 588222 203994
rect 588458 203758 588542 203994
rect 588778 203758 588810 203994
rect 588190 167994 588810 203758
rect 588190 167758 588222 167994
rect 588458 167758 588542 167994
rect 588778 167758 588810 167994
rect 588190 131994 588810 167758
rect 588190 131758 588222 131994
rect 588458 131758 588542 131994
rect 588778 131758 588810 131994
rect 588190 95994 588810 131758
rect 588190 95758 588222 95994
rect 588458 95758 588542 95994
rect 588778 95758 588810 95994
rect 588190 59994 588810 95758
rect 588190 59758 588222 59994
rect 588458 59758 588542 59994
rect 588778 59758 588810 59994
rect 588190 23994 588810 59758
rect 588190 23758 588222 23994
rect 588458 23758 588542 23994
rect 588778 23758 588810 23994
rect 588190 -3226 588810 23758
rect 588190 -3462 588222 -3226
rect 588458 -3462 588542 -3226
rect 588778 -3462 588810 -3226
rect 588190 -3546 588810 -3462
rect 588190 -3782 588222 -3546
rect 588458 -3782 588542 -3546
rect 588778 -3782 588810 -3546
rect 588190 -3814 588810 -3782
rect 589150 693694 589770 708122
rect 589150 693458 589182 693694
rect 589418 693458 589502 693694
rect 589738 693458 589770 693694
rect 589150 657694 589770 693458
rect 589150 657458 589182 657694
rect 589418 657458 589502 657694
rect 589738 657458 589770 657694
rect 589150 621694 589770 657458
rect 589150 621458 589182 621694
rect 589418 621458 589502 621694
rect 589738 621458 589770 621694
rect 589150 585694 589770 621458
rect 589150 585458 589182 585694
rect 589418 585458 589502 585694
rect 589738 585458 589770 585694
rect 589150 549694 589770 585458
rect 589150 549458 589182 549694
rect 589418 549458 589502 549694
rect 589738 549458 589770 549694
rect 589150 513694 589770 549458
rect 589150 513458 589182 513694
rect 589418 513458 589502 513694
rect 589738 513458 589770 513694
rect 589150 477694 589770 513458
rect 589150 477458 589182 477694
rect 589418 477458 589502 477694
rect 589738 477458 589770 477694
rect 589150 441694 589770 477458
rect 589150 441458 589182 441694
rect 589418 441458 589502 441694
rect 589738 441458 589770 441694
rect 589150 405694 589770 441458
rect 589150 405458 589182 405694
rect 589418 405458 589502 405694
rect 589738 405458 589770 405694
rect 589150 369694 589770 405458
rect 589150 369458 589182 369694
rect 589418 369458 589502 369694
rect 589738 369458 589770 369694
rect 589150 333694 589770 369458
rect 589150 333458 589182 333694
rect 589418 333458 589502 333694
rect 589738 333458 589770 333694
rect 589150 297694 589770 333458
rect 589150 297458 589182 297694
rect 589418 297458 589502 297694
rect 589738 297458 589770 297694
rect 589150 261694 589770 297458
rect 589150 261458 589182 261694
rect 589418 261458 589502 261694
rect 589738 261458 589770 261694
rect 589150 225694 589770 261458
rect 589150 225458 589182 225694
rect 589418 225458 589502 225694
rect 589738 225458 589770 225694
rect 589150 189694 589770 225458
rect 589150 189458 589182 189694
rect 589418 189458 589502 189694
rect 589738 189458 589770 189694
rect 589150 153694 589770 189458
rect 589150 153458 589182 153694
rect 589418 153458 589502 153694
rect 589738 153458 589770 153694
rect 589150 117694 589770 153458
rect 589150 117458 589182 117694
rect 589418 117458 589502 117694
rect 589738 117458 589770 117694
rect 589150 81694 589770 117458
rect 589150 81458 589182 81694
rect 589418 81458 589502 81694
rect 589738 81458 589770 81694
rect 589150 45694 589770 81458
rect 589150 45458 589182 45694
rect 589418 45458 589502 45694
rect 589738 45458 589770 45694
rect 589150 9694 589770 45458
rect 589150 9458 589182 9694
rect 589418 9458 589502 9694
rect 589738 9458 589770 9694
rect 589150 -4186 589770 9458
rect 589150 -4422 589182 -4186
rect 589418 -4422 589502 -4186
rect 589738 -4422 589770 -4186
rect 589150 -4506 589770 -4422
rect 589150 -4742 589182 -4506
rect 589418 -4742 589502 -4506
rect 589738 -4742 589770 -4506
rect 589150 -4774 589770 -4742
rect 590110 675694 590730 709082
rect 590110 675458 590142 675694
rect 590378 675458 590462 675694
rect 590698 675458 590730 675694
rect 590110 639694 590730 675458
rect 590110 639458 590142 639694
rect 590378 639458 590462 639694
rect 590698 639458 590730 639694
rect 590110 603694 590730 639458
rect 590110 603458 590142 603694
rect 590378 603458 590462 603694
rect 590698 603458 590730 603694
rect 590110 567694 590730 603458
rect 590110 567458 590142 567694
rect 590378 567458 590462 567694
rect 590698 567458 590730 567694
rect 590110 531694 590730 567458
rect 590110 531458 590142 531694
rect 590378 531458 590462 531694
rect 590698 531458 590730 531694
rect 590110 495694 590730 531458
rect 590110 495458 590142 495694
rect 590378 495458 590462 495694
rect 590698 495458 590730 495694
rect 590110 459694 590730 495458
rect 590110 459458 590142 459694
rect 590378 459458 590462 459694
rect 590698 459458 590730 459694
rect 590110 423694 590730 459458
rect 590110 423458 590142 423694
rect 590378 423458 590462 423694
rect 590698 423458 590730 423694
rect 590110 387694 590730 423458
rect 590110 387458 590142 387694
rect 590378 387458 590462 387694
rect 590698 387458 590730 387694
rect 590110 351694 590730 387458
rect 590110 351458 590142 351694
rect 590378 351458 590462 351694
rect 590698 351458 590730 351694
rect 590110 315694 590730 351458
rect 590110 315458 590142 315694
rect 590378 315458 590462 315694
rect 590698 315458 590730 315694
rect 590110 279694 590730 315458
rect 590110 279458 590142 279694
rect 590378 279458 590462 279694
rect 590698 279458 590730 279694
rect 590110 243694 590730 279458
rect 590110 243458 590142 243694
rect 590378 243458 590462 243694
rect 590698 243458 590730 243694
rect 590110 207694 590730 243458
rect 590110 207458 590142 207694
rect 590378 207458 590462 207694
rect 590698 207458 590730 207694
rect 590110 171694 590730 207458
rect 590110 171458 590142 171694
rect 590378 171458 590462 171694
rect 590698 171458 590730 171694
rect 590110 135694 590730 171458
rect 590110 135458 590142 135694
rect 590378 135458 590462 135694
rect 590698 135458 590730 135694
rect 590110 99694 590730 135458
rect 590110 99458 590142 99694
rect 590378 99458 590462 99694
rect 590698 99458 590730 99694
rect 590110 63694 590730 99458
rect 590110 63458 590142 63694
rect 590378 63458 590462 63694
rect 590698 63458 590730 63694
rect 590110 27694 590730 63458
rect 590110 27458 590142 27694
rect 590378 27458 590462 27694
rect 590698 27458 590730 27694
rect 590110 -5146 590730 27458
rect 590110 -5382 590142 -5146
rect 590378 -5382 590462 -5146
rect 590698 -5382 590730 -5146
rect 590110 -5466 590730 -5382
rect 590110 -5702 590142 -5466
rect 590378 -5702 590462 -5466
rect 590698 -5702 590730 -5466
rect 590110 -5734 590730 -5702
rect 591070 697394 591690 710042
rect 591070 697158 591102 697394
rect 591338 697158 591422 697394
rect 591658 697158 591690 697394
rect 591070 661394 591690 697158
rect 591070 661158 591102 661394
rect 591338 661158 591422 661394
rect 591658 661158 591690 661394
rect 591070 625394 591690 661158
rect 591070 625158 591102 625394
rect 591338 625158 591422 625394
rect 591658 625158 591690 625394
rect 591070 589394 591690 625158
rect 591070 589158 591102 589394
rect 591338 589158 591422 589394
rect 591658 589158 591690 589394
rect 591070 553394 591690 589158
rect 591070 553158 591102 553394
rect 591338 553158 591422 553394
rect 591658 553158 591690 553394
rect 591070 517394 591690 553158
rect 591070 517158 591102 517394
rect 591338 517158 591422 517394
rect 591658 517158 591690 517394
rect 591070 481394 591690 517158
rect 591070 481158 591102 481394
rect 591338 481158 591422 481394
rect 591658 481158 591690 481394
rect 591070 445394 591690 481158
rect 591070 445158 591102 445394
rect 591338 445158 591422 445394
rect 591658 445158 591690 445394
rect 591070 409394 591690 445158
rect 591070 409158 591102 409394
rect 591338 409158 591422 409394
rect 591658 409158 591690 409394
rect 591070 373394 591690 409158
rect 591070 373158 591102 373394
rect 591338 373158 591422 373394
rect 591658 373158 591690 373394
rect 591070 337394 591690 373158
rect 591070 337158 591102 337394
rect 591338 337158 591422 337394
rect 591658 337158 591690 337394
rect 591070 301394 591690 337158
rect 591070 301158 591102 301394
rect 591338 301158 591422 301394
rect 591658 301158 591690 301394
rect 591070 265394 591690 301158
rect 591070 265158 591102 265394
rect 591338 265158 591422 265394
rect 591658 265158 591690 265394
rect 591070 229394 591690 265158
rect 591070 229158 591102 229394
rect 591338 229158 591422 229394
rect 591658 229158 591690 229394
rect 591070 193394 591690 229158
rect 591070 193158 591102 193394
rect 591338 193158 591422 193394
rect 591658 193158 591690 193394
rect 591070 157394 591690 193158
rect 591070 157158 591102 157394
rect 591338 157158 591422 157394
rect 591658 157158 591690 157394
rect 591070 121394 591690 157158
rect 591070 121158 591102 121394
rect 591338 121158 591422 121394
rect 591658 121158 591690 121394
rect 591070 85394 591690 121158
rect 591070 85158 591102 85394
rect 591338 85158 591422 85394
rect 591658 85158 591690 85394
rect 591070 49394 591690 85158
rect 591070 49158 591102 49394
rect 591338 49158 591422 49394
rect 591658 49158 591690 49394
rect 591070 13394 591690 49158
rect 591070 13158 591102 13394
rect 591338 13158 591422 13394
rect 591658 13158 591690 13394
rect 591070 -6106 591690 13158
rect 591070 -6342 591102 -6106
rect 591338 -6342 591422 -6106
rect 591658 -6342 591690 -6106
rect 591070 -6426 591690 -6342
rect 591070 -6662 591102 -6426
rect 591338 -6662 591422 -6426
rect 591658 -6662 591690 -6426
rect 591070 -6694 591690 -6662
rect 592030 679394 592650 711002
rect 592030 679158 592062 679394
rect 592298 679158 592382 679394
rect 592618 679158 592650 679394
rect 592030 643394 592650 679158
rect 592030 643158 592062 643394
rect 592298 643158 592382 643394
rect 592618 643158 592650 643394
rect 592030 607394 592650 643158
rect 592030 607158 592062 607394
rect 592298 607158 592382 607394
rect 592618 607158 592650 607394
rect 592030 571394 592650 607158
rect 592030 571158 592062 571394
rect 592298 571158 592382 571394
rect 592618 571158 592650 571394
rect 592030 535394 592650 571158
rect 592030 535158 592062 535394
rect 592298 535158 592382 535394
rect 592618 535158 592650 535394
rect 592030 499394 592650 535158
rect 592030 499158 592062 499394
rect 592298 499158 592382 499394
rect 592618 499158 592650 499394
rect 592030 463394 592650 499158
rect 592030 463158 592062 463394
rect 592298 463158 592382 463394
rect 592618 463158 592650 463394
rect 592030 427394 592650 463158
rect 592030 427158 592062 427394
rect 592298 427158 592382 427394
rect 592618 427158 592650 427394
rect 592030 391394 592650 427158
rect 592030 391158 592062 391394
rect 592298 391158 592382 391394
rect 592618 391158 592650 391394
rect 592030 355394 592650 391158
rect 592030 355158 592062 355394
rect 592298 355158 592382 355394
rect 592618 355158 592650 355394
rect 592030 319394 592650 355158
rect 592030 319158 592062 319394
rect 592298 319158 592382 319394
rect 592618 319158 592650 319394
rect 592030 283394 592650 319158
rect 592030 283158 592062 283394
rect 592298 283158 592382 283394
rect 592618 283158 592650 283394
rect 592030 247394 592650 283158
rect 592030 247158 592062 247394
rect 592298 247158 592382 247394
rect 592618 247158 592650 247394
rect 592030 211394 592650 247158
rect 592030 211158 592062 211394
rect 592298 211158 592382 211394
rect 592618 211158 592650 211394
rect 592030 175394 592650 211158
rect 592030 175158 592062 175394
rect 592298 175158 592382 175394
rect 592618 175158 592650 175394
rect 592030 139394 592650 175158
rect 592030 139158 592062 139394
rect 592298 139158 592382 139394
rect 592618 139158 592650 139394
rect 592030 103394 592650 139158
rect 592030 103158 592062 103394
rect 592298 103158 592382 103394
rect 592618 103158 592650 103394
rect 592030 67394 592650 103158
rect 592030 67158 592062 67394
rect 592298 67158 592382 67394
rect 592618 67158 592650 67394
rect 592030 31394 592650 67158
rect 592030 31158 592062 31394
rect 592298 31158 592382 31394
rect 592618 31158 592650 31394
rect 569904 -7302 570086 -7066
rect 570322 -7302 570504 -7066
rect 569904 -7386 570504 -7302
rect 569904 -7622 570086 -7386
rect 570322 -7622 570504 -7386
rect 569904 -7654 570504 -7622
rect 592030 -7066 592650 31158
rect 592030 -7302 592062 -7066
rect 592298 -7302 592382 -7066
rect 592618 -7302 592650 -7066
rect 592030 -7386 592650 -7302
rect 592030 -7622 592062 -7386
rect 592298 -7622 592382 -7386
rect 592618 -7622 592650 -7386
rect 592030 -7654 592650 -7622
<< via4 >>
rect -8694 711322 -8458 711558
rect -8374 711322 -8138 711558
rect -8694 711002 -8458 711238
rect -8374 711002 -8138 711238
rect -8694 679158 -8458 679394
rect -8374 679158 -8138 679394
rect -8694 643158 -8458 643394
rect -8374 643158 -8138 643394
rect -8694 607158 -8458 607394
rect -8374 607158 -8138 607394
rect -8694 571158 -8458 571394
rect -8374 571158 -8138 571394
rect -8694 535158 -8458 535394
rect -8374 535158 -8138 535394
rect -8694 499158 -8458 499394
rect -8374 499158 -8138 499394
rect -8694 463158 -8458 463394
rect -8374 463158 -8138 463394
rect -8694 427158 -8458 427394
rect -8374 427158 -8138 427394
rect -8694 391158 -8458 391394
rect -8374 391158 -8138 391394
rect -8694 355158 -8458 355394
rect -8374 355158 -8138 355394
rect -8694 319158 -8458 319394
rect -8374 319158 -8138 319394
rect -8694 283158 -8458 283394
rect -8374 283158 -8138 283394
rect -8694 247158 -8458 247394
rect -8374 247158 -8138 247394
rect -8694 211158 -8458 211394
rect -8374 211158 -8138 211394
rect -8694 175158 -8458 175394
rect -8374 175158 -8138 175394
rect -8694 139158 -8458 139394
rect -8374 139158 -8138 139394
rect -8694 103158 -8458 103394
rect -8374 103158 -8138 103394
rect -8694 67158 -8458 67394
rect -8374 67158 -8138 67394
rect -8694 31158 -8458 31394
rect -8374 31158 -8138 31394
rect -7734 710362 -7498 710598
rect -7414 710362 -7178 710598
rect -7734 710042 -7498 710278
rect -7414 710042 -7178 710278
rect 12086 710362 12322 710598
rect 12086 710042 12322 710278
rect -7734 697158 -7498 697394
rect -7414 697158 -7178 697394
rect -7734 661158 -7498 661394
rect -7414 661158 -7178 661394
rect -7734 625158 -7498 625394
rect -7414 625158 -7178 625394
rect -7734 589158 -7498 589394
rect -7414 589158 -7178 589394
rect -7734 553158 -7498 553394
rect -7414 553158 -7178 553394
rect -7734 517158 -7498 517394
rect -7414 517158 -7178 517394
rect -7734 481158 -7498 481394
rect -7414 481158 -7178 481394
rect -7734 445158 -7498 445394
rect -7414 445158 -7178 445394
rect -7734 409158 -7498 409394
rect -7414 409158 -7178 409394
rect -7734 373158 -7498 373394
rect -7414 373158 -7178 373394
rect -7734 337158 -7498 337394
rect -7414 337158 -7178 337394
rect -7734 301158 -7498 301394
rect -7414 301158 -7178 301394
rect -7734 265158 -7498 265394
rect -7414 265158 -7178 265394
rect -7734 229158 -7498 229394
rect -7414 229158 -7178 229394
rect -7734 193158 -7498 193394
rect -7414 193158 -7178 193394
rect -7734 157158 -7498 157394
rect -7414 157158 -7178 157394
rect -7734 121158 -7498 121394
rect -7414 121158 -7178 121394
rect -7734 85158 -7498 85394
rect -7414 85158 -7178 85394
rect -7734 49158 -7498 49394
rect -7414 49158 -7178 49394
rect -7734 13158 -7498 13394
rect -7414 13158 -7178 13394
rect -6774 709402 -6538 709638
rect -6454 709402 -6218 709638
rect -6774 709082 -6538 709318
rect -6454 709082 -6218 709318
rect -6774 675458 -6538 675694
rect -6454 675458 -6218 675694
rect -6774 639458 -6538 639694
rect -6454 639458 -6218 639694
rect -6774 603458 -6538 603694
rect -6454 603458 -6218 603694
rect -6774 567458 -6538 567694
rect -6454 567458 -6218 567694
rect -6774 531458 -6538 531694
rect -6454 531458 -6218 531694
rect -6774 495458 -6538 495694
rect -6454 495458 -6218 495694
rect -6774 459458 -6538 459694
rect -6454 459458 -6218 459694
rect -6774 423458 -6538 423694
rect -6454 423458 -6218 423694
rect -6774 387458 -6538 387694
rect -6454 387458 -6218 387694
rect -6774 351458 -6538 351694
rect -6454 351458 -6218 351694
rect -6774 315458 -6538 315694
rect -6454 315458 -6218 315694
rect -6774 279458 -6538 279694
rect -6454 279458 -6218 279694
rect -6774 243458 -6538 243694
rect -6454 243458 -6218 243694
rect -6774 207458 -6538 207694
rect -6454 207458 -6218 207694
rect -6774 171458 -6538 171694
rect -6454 171458 -6218 171694
rect -6774 135458 -6538 135694
rect -6454 135458 -6218 135694
rect -6774 99458 -6538 99694
rect -6454 99458 -6218 99694
rect -6774 63458 -6538 63694
rect -6454 63458 -6218 63694
rect -6774 27458 -6538 27694
rect -6454 27458 -6218 27694
rect -5814 708442 -5578 708678
rect -5494 708442 -5258 708678
rect -5814 708122 -5578 708358
rect -5494 708122 -5258 708358
rect 8386 708442 8622 708678
rect 8386 708122 8622 708358
rect -5814 693458 -5578 693694
rect -5494 693458 -5258 693694
rect -5814 657458 -5578 657694
rect -5494 657458 -5258 657694
rect -5814 621458 -5578 621694
rect -5494 621458 -5258 621694
rect -5814 585458 -5578 585694
rect -5494 585458 -5258 585694
rect -5814 549458 -5578 549694
rect -5494 549458 -5258 549694
rect -5814 513458 -5578 513694
rect -5494 513458 -5258 513694
rect -5814 477458 -5578 477694
rect -5494 477458 -5258 477694
rect -5814 441458 -5578 441694
rect -5494 441458 -5258 441694
rect -5814 405458 -5578 405694
rect -5494 405458 -5258 405694
rect -5814 369458 -5578 369694
rect -5494 369458 -5258 369694
rect -5814 333458 -5578 333694
rect -5494 333458 -5258 333694
rect -5814 297458 -5578 297694
rect -5494 297458 -5258 297694
rect -5814 261458 -5578 261694
rect -5494 261458 -5258 261694
rect -5814 225458 -5578 225694
rect -5494 225458 -5258 225694
rect -5814 189458 -5578 189694
rect -5494 189458 -5258 189694
rect -5814 153458 -5578 153694
rect -5494 153458 -5258 153694
rect -5814 117458 -5578 117694
rect -5494 117458 -5258 117694
rect -5814 81458 -5578 81694
rect -5494 81458 -5258 81694
rect -5814 45458 -5578 45694
rect -5494 45458 -5258 45694
rect -5814 9458 -5578 9694
rect -5494 9458 -5258 9694
rect -4854 707482 -4618 707718
rect -4534 707482 -4298 707718
rect -4854 707162 -4618 707398
rect -4534 707162 -4298 707398
rect -4854 671758 -4618 671994
rect -4534 671758 -4298 671994
rect -4854 635758 -4618 635994
rect -4534 635758 -4298 635994
rect -4854 599758 -4618 599994
rect -4534 599758 -4298 599994
rect -4854 563758 -4618 563994
rect -4534 563758 -4298 563994
rect -4854 527758 -4618 527994
rect -4534 527758 -4298 527994
rect -4854 491758 -4618 491994
rect -4534 491758 -4298 491994
rect -4854 455758 -4618 455994
rect -4534 455758 -4298 455994
rect -4854 419758 -4618 419994
rect -4534 419758 -4298 419994
rect -4854 383758 -4618 383994
rect -4534 383758 -4298 383994
rect -4854 347758 -4618 347994
rect -4534 347758 -4298 347994
rect -4854 311758 -4618 311994
rect -4534 311758 -4298 311994
rect -4854 275758 -4618 275994
rect -4534 275758 -4298 275994
rect -4854 239758 -4618 239994
rect -4534 239758 -4298 239994
rect -4854 203758 -4618 203994
rect -4534 203758 -4298 203994
rect -4854 167758 -4618 167994
rect -4534 167758 -4298 167994
rect -4854 131758 -4618 131994
rect -4534 131758 -4298 131994
rect -4854 95758 -4618 95994
rect -4534 95758 -4298 95994
rect -4854 59758 -4618 59994
rect -4534 59758 -4298 59994
rect -4854 23758 -4618 23994
rect -4534 23758 -4298 23994
rect -3894 706522 -3658 706758
rect -3574 706522 -3338 706758
rect -3894 706202 -3658 706438
rect -3574 706202 -3338 706438
rect 4686 706522 4922 706758
rect 4686 706202 4922 706438
rect -3894 689758 -3658 689994
rect -3574 689758 -3338 689994
rect -3894 653758 -3658 653994
rect -3574 653758 -3338 653994
rect -3894 617758 -3658 617994
rect -3574 617758 -3338 617994
rect -3894 581758 -3658 581994
rect -3574 581758 -3338 581994
rect -3894 545758 -3658 545994
rect -3574 545758 -3338 545994
rect -3894 509758 -3658 509994
rect -3574 509758 -3338 509994
rect -3894 473758 -3658 473994
rect -3574 473758 -3338 473994
rect -3894 437758 -3658 437994
rect -3574 437758 -3338 437994
rect -3894 401758 -3658 401994
rect -3574 401758 -3338 401994
rect -3894 365758 -3658 365994
rect -3574 365758 -3338 365994
rect -3894 329758 -3658 329994
rect -3574 329758 -3338 329994
rect -3894 293758 -3658 293994
rect -3574 293758 -3338 293994
rect -3894 257758 -3658 257994
rect -3574 257758 -3338 257994
rect -3894 221758 -3658 221994
rect -3574 221758 -3338 221994
rect -3894 185758 -3658 185994
rect -3574 185758 -3338 185994
rect -3894 149758 -3658 149994
rect -3574 149758 -3338 149994
rect -3894 113758 -3658 113994
rect -3574 113758 -3338 113994
rect -3894 77758 -3658 77994
rect -3574 77758 -3338 77994
rect -3894 41758 -3658 41994
rect -3574 41758 -3338 41994
rect -3894 5758 -3658 5994
rect -3574 5758 -3338 5994
rect -2934 705562 -2698 705798
rect -2614 705562 -2378 705798
rect -2934 705242 -2698 705478
rect -2614 705242 -2378 705478
rect -2934 668058 -2698 668294
rect -2614 668058 -2378 668294
rect -2934 632058 -2698 632294
rect -2614 632058 -2378 632294
rect -2934 596058 -2698 596294
rect -2614 596058 -2378 596294
rect -2934 560058 -2698 560294
rect -2614 560058 -2378 560294
rect -2934 524058 -2698 524294
rect -2614 524058 -2378 524294
rect -2934 488058 -2698 488294
rect -2614 488058 -2378 488294
rect -2934 452058 -2698 452294
rect -2614 452058 -2378 452294
rect -2934 416058 -2698 416294
rect -2614 416058 -2378 416294
rect -2934 380058 -2698 380294
rect -2614 380058 -2378 380294
rect -2934 344058 -2698 344294
rect -2614 344058 -2378 344294
rect -2934 308058 -2698 308294
rect -2614 308058 -2378 308294
rect -2934 272058 -2698 272294
rect -2614 272058 -2378 272294
rect -2934 236058 -2698 236294
rect -2614 236058 -2378 236294
rect -2934 200058 -2698 200294
rect -2614 200058 -2378 200294
rect -2934 164058 -2698 164294
rect -2614 164058 -2378 164294
rect -2934 128058 -2698 128294
rect -2614 128058 -2378 128294
rect -2934 92058 -2698 92294
rect -2614 92058 -2378 92294
rect -2934 56058 -2698 56294
rect -2614 56058 -2378 56294
rect -2934 20058 -2698 20294
rect -2614 20058 -2378 20294
rect -1974 704602 -1738 704838
rect -1654 704602 -1418 704838
rect -1974 704282 -1738 704518
rect -1654 704282 -1418 704518
rect -1974 686058 -1738 686294
rect -1654 686058 -1418 686294
rect -1974 650058 -1738 650294
rect -1654 650058 -1418 650294
rect -1974 614058 -1738 614294
rect -1654 614058 -1418 614294
rect -1974 578058 -1738 578294
rect -1654 578058 -1418 578294
rect -1974 542058 -1738 542294
rect -1654 542058 -1418 542294
rect -1974 506058 -1738 506294
rect -1654 506058 -1418 506294
rect -1974 470058 -1738 470294
rect -1654 470058 -1418 470294
rect -1974 434058 -1738 434294
rect -1654 434058 -1418 434294
rect -1974 398058 -1738 398294
rect -1654 398058 -1418 398294
rect -1974 362058 -1738 362294
rect -1654 362058 -1418 362294
rect -1974 326058 -1738 326294
rect -1654 326058 -1418 326294
rect -1974 290058 -1738 290294
rect -1654 290058 -1418 290294
rect -1974 254058 -1738 254294
rect -1654 254058 -1418 254294
rect -1974 218058 -1738 218294
rect -1654 218058 -1418 218294
rect -1974 182058 -1738 182294
rect -1654 182058 -1418 182294
rect -1974 146058 -1738 146294
rect -1654 146058 -1418 146294
rect -1974 110058 -1738 110294
rect -1654 110058 -1418 110294
rect -1974 74058 -1738 74294
rect -1654 74058 -1418 74294
rect -1974 38058 -1738 38294
rect -1654 38058 -1418 38294
rect -1974 2058 -1738 2294
rect -1654 2058 -1418 2294
rect -1974 -582 -1738 -346
rect -1654 -582 -1418 -346
rect -1974 -902 -1738 -666
rect -1654 -902 -1418 -666
rect 986 704602 1222 704838
rect 986 704282 1222 704518
rect 986 686058 1222 686294
rect 986 650058 1222 650294
rect 986 614058 1222 614294
rect 986 578058 1222 578294
rect 986 542058 1222 542294
rect 986 506058 1222 506294
rect 986 470058 1222 470294
rect 986 434058 1222 434294
rect 986 398058 1222 398294
rect 986 362058 1222 362294
rect 986 326058 1222 326294
rect 986 290058 1222 290294
rect 986 254058 1222 254294
rect 986 218058 1222 218294
rect 986 182058 1222 182294
rect 986 146058 1222 146294
rect 986 110058 1222 110294
rect 986 74058 1222 74294
rect 986 38058 1222 38294
rect 986 2058 1222 2294
rect 986 -582 1222 -346
rect 986 -902 1222 -666
rect -2934 -1542 -2698 -1306
rect -2614 -1542 -2378 -1306
rect -2934 -1862 -2698 -1626
rect -2614 -1862 -2378 -1626
rect 4686 689758 4922 689994
rect 4686 653758 4922 653994
rect 4686 617758 4922 617994
rect 4686 581758 4922 581994
rect 4686 545758 4922 545994
rect 4686 509758 4922 509994
rect 4686 473758 4922 473994
rect 4686 437758 4922 437994
rect 4686 401758 4922 401994
rect 4686 365758 4922 365994
rect 4686 329758 4922 329994
rect 4686 293758 4922 293994
rect 4686 257758 4922 257994
rect 4686 221758 4922 221994
rect 4686 185758 4922 185994
rect 4686 149758 4922 149994
rect 4686 113758 4922 113994
rect 4686 77758 4922 77994
rect 4686 41758 4922 41994
rect 4686 5758 4922 5994
rect -3894 -2502 -3658 -2266
rect -3574 -2502 -3338 -2266
rect -3894 -2822 -3658 -2586
rect -3574 -2822 -3338 -2586
rect 4686 -2502 4922 -2266
rect 4686 -2822 4922 -2586
rect -4854 -3462 -4618 -3226
rect -4534 -3462 -4298 -3226
rect -4854 -3782 -4618 -3546
rect -4534 -3782 -4298 -3546
rect 8386 693458 8622 693694
rect 8386 657458 8622 657694
rect 8386 621458 8622 621694
rect 8386 585458 8622 585694
rect 8386 549458 8622 549694
rect 8386 513458 8622 513694
rect 8386 477458 8622 477694
rect 8386 441458 8622 441694
rect 8386 405458 8622 405694
rect 8386 369458 8622 369694
rect 8386 333458 8622 333694
rect 8386 297458 8622 297694
rect 8386 261458 8622 261694
rect 8386 225458 8622 225694
rect 8386 189458 8622 189694
rect 8386 153458 8622 153694
rect 8386 117458 8622 117694
rect 8386 81458 8622 81694
rect 8386 45458 8622 45694
rect 8386 9458 8622 9694
rect -5814 -4422 -5578 -4186
rect -5494 -4422 -5258 -4186
rect -5814 -4742 -5578 -4506
rect -5494 -4742 -5258 -4506
rect 8386 -4422 8622 -4186
rect 8386 -4742 8622 -4506
rect -6774 -5382 -6538 -5146
rect -6454 -5382 -6218 -5146
rect -6774 -5702 -6538 -5466
rect -6454 -5702 -6218 -5466
rect 30086 711322 30322 711558
rect 30086 711002 30322 711238
rect 26386 709402 26622 709638
rect 26386 709082 26622 709318
rect 22686 707482 22922 707718
rect 22686 707162 22922 707398
rect 12086 697158 12322 697394
rect 12086 661158 12322 661394
rect 12086 625158 12322 625394
rect 12086 589158 12322 589394
rect 12086 553158 12322 553394
rect 12086 517158 12322 517394
rect 12086 481158 12322 481394
rect 12086 445158 12322 445394
rect 12086 409158 12322 409394
rect 12086 373158 12322 373394
rect 12086 337158 12322 337394
rect 12086 301158 12322 301394
rect 12086 265158 12322 265394
rect 12086 229158 12322 229394
rect 12086 193158 12322 193394
rect 12086 157158 12322 157394
rect 12086 121158 12322 121394
rect 12086 85158 12322 85394
rect 12086 49158 12322 49394
rect 12086 13158 12322 13394
rect -7734 -6342 -7498 -6106
rect -7414 -6342 -7178 -6106
rect -7734 -6662 -7498 -6426
rect -7414 -6662 -7178 -6426
rect 18986 705562 19222 705798
rect 18986 705242 19222 705478
rect 18986 668058 19222 668294
rect 18986 632058 19222 632294
rect 18986 596058 19222 596294
rect 18986 560058 19222 560294
rect 18986 524058 19222 524294
rect 18986 488058 19222 488294
rect 18986 452058 19222 452294
rect 18986 416058 19222 416294
rect 18986 380058 19222 380294
rect 18986 344058 19222 344294
rect 18986 308058 19222 308294
rect 18986 272058 19222 272294
rect 18986 236058 19222 236294
rect 18986 200058 19222 200294
rect 18986 164058 19222 164294
rect 18986 128058 19222 128294
rect 18986 92058 19222 92294
rect 18986 56058 19222 56294
rect 18986 20058 19222 20294
rect 18986 -1542 19222 -1306
rect 18986 -1862 19222 -1626
rect 22686 671758 22922 671994
rect 22686 635758 22922 635994
rect 22686 599758 22922 599994
rect 22686 563758 22922 563994
rect 22686 527758 22922 527994
rect 22686 491758 22922 491994
rect 22686 455758 22922 455994
rect 22686 419758 22922 419994
rect 22686 383758 22922 383994
rect 22686 347758 22922 347994
rect 22686 311758 22922 311994
rect 22686 275758 22922 275994
rect 22686 239758 22922 239994
rect 22686 203758 22922 203994
rect 22686 167758 22922 167994
rect 22686 131758 22922 131994
rect 22686 95758 22922 95994
rect 22686 59758 22922 59994
rect 22686 23758 22922 23994
rect 22686 -3462 22922 -3226
rect 22686 -3782 22922 -3546
rect 26386 675458 26622 675694
rect 26386 639458 26622 639694
rect 26386 603458 26622 603694
rect 26386 567458 26622 567694
rect 26386 531458 26622 531694
rect 26386 495458 26622 495694
rect 26386 459458 26622 459694
rect 26386 423458 26622 423694
rect 26386 387458 26622 387694
rect 26386 351458 26622 351694
rect 26386 315458 26622 315694
rect 26386 279458 26622 279694
rect 26386 243458 26622 243694
rect 26386 207458 26622 207694
rect 26386 171458 26622 171694
rect 26386 135458 26622 135694
rect 26386 99458 26622 99694
rect 26386 63458 26622 63694
rect 26386 27458 26622 27694
rect 26386 -5382 26622 -5146
rect 26386 -5702 26622 -5466
rect 48086 710362 48322 710598
rect 48086 710042 48322 710278
rect 44386 708442 44622 708678
rect 44386 708122 44622 708358
rect 40686 706522 40922 706758
rect 40686 706202 40922 706438
rect 30086 679158 30322 679394
rect 30086 643158 30322 643394
rect 30086 607158 30322 607394
rect 30086 571158 30322 571394
rect 30086 535158 30322 535394
rect 30086 499158 30322 499394
rect 30086 463158 30322 463394
rect 30086 427158 30322 427394
rect 30086 391158 30322 391394
rect 30086 355158 30322 355394
rect 30086 319158 30322 319394
rect 30086 283158 30322 283394
rect 30086 247158 30322 247394
rect 30086 211158 30322 211394
rect 30086 175158 30322 175394
rect 30086 139158 30322 139394
rect 30086 103158 30322 103394
rect 30086 67158 30322 67394
rect 30086 31158 30322 31394
rect 12086 -6342 12322 -6106
rect 12086 -6662 12322 -6426
rect -8694 -7302 -8458 -7066
rect -8374 -7302 -8138 -7066
rect -8694 -7622 -8458 -7386
rect -8374 -7622 -8138 -7386
rect 36986 704602 37222 704838
rect 36986 704282 37222 704518
rect 36986 686058 37222 686294
rect 36986 650058 37222 650294
rect 36986 614058 37222 614294
rect 36986 578058 37222 578294
rect 36986 542058 37222 542294
rect 36986 506058 37222 506294
rect 36986 470058 37222 470294
rect 36986 434058 37222 434294
rect 40686 689758 40922 689994
rect 40686 653758 40922 653994
rect 40686 617758 40922 617994
rect 40686 581758 40922 581994
rect 40686 545758 40922 545994
rect 40686 509758 40922 509994
rect 40686 473758 40922 473994
rect 40686 437758 40922 437994
rect 44386 693458 44622 693694
rect 44386 657458 44622 657694
rect 44386 621458 44622 621694
rect 44386 585458 44622 585694
rect 44386 549458 44622 549694
rect 44386 513458 44622 513694
rect 44386 477458 44622 477694
rect 44386 441458 44622 441694
rect 66086 711322 66322 711558
rect 66086 711002 66322 711238
rect 62386 709402 62622 709638
rect 62386 709082 62622 709318
rect 58686 707482 58922 707718
rect 58686 707162 58922 707398
rect 48086 697158 48322 697394
rect 48086 661158 48322 661394
rect 48086 625158 48322 625394
rect 48086 589158 48322 589394
rect 48086 553158 48322 553394
rect 48086 517158 48322 517394
rect 48086 481158 48322 481394
rect 48086 445158 48322 445394
rect 54986 705562 55222 705798
rect 54986 705242 55222 705478
rect 54986 668058 55222 668294
rect 54986 632058 55222 632294
rect 54986 596058 55222 596294
rect 54986 560058 55222 560294
rect 54986 524058 55222 524294
rect 54986 488058 55222 488294
rect 54986 452058 55222 452294
rect 58686 671758 58922 671994
rect 58686 635758 58922 635994
rect 58686 599758 58922 599994
rect 58686 563758 58922 563994
rect 58686 527758 58922 527994
rect 58686 491758 58922 491994
rect 58686 455758 58922 455994
rect 62386 675458 62622 675694
rect 62386 639458 62622 639694
rect 62386 603458 62622 603694
rect 62386 567458 62622 567694
rect 62386 531458 62622 531694
rect 62386 495458 62622 495694
rect 62386 459458 62622 459694
rect 84086 710362 84322 710598
rect 84086 710042 84322 710278
rect 80386 708442 80622 708678
rect 80386 708122 80622 708358
rect 76686 706522 76922 706758
rect 76686 706202 76922 706438
rect 66086 679158 66322 679394
rect 66086 643158 66322 643394
rect 66086 607158 66322 607394
rect 66086 571158 66322 571394
rect 66086 535158 66322 535394
rect 66086 499158 66322 499394
rect 66086 463158 66322 463394
rect 66086 427158 66322 427394
rect 72986 704602 73222 704838
rect 72986 704282 73222 704518
rect 72986 686058 73222 686294
rect 72986 650058 73222 650294
rect 72986 614058 73222 614294
rect 72986 578058 73222 578294
rect 72986 542058 73222 542294
rect 72986 506058 73222 506294
rect 72986 470058 73222 470294
rect 72986 434058 73222 434294
rect 76686 689758 76922 689994
rect 76686 653758 76922 653994
rect 76686 617758 76922 617994
rect 76686 581758 76922 581994
rect 76686 545758 76922 545994
rect 76686 509758 76922 509994
rect 76686 473758 76922 473994
rect 76686 437758 76922 437994
rect 80386 693458 80622 693694
rect 80386 657458 80622 657694
rect 80386 621458 80622 621694
rect 80386 585458 80622 585694
rect 80386 549458 80622 549694
rect 80386 513458 80622 513694
rect 80386 477458 80622 477694
rect 80386 441458 80622 441694
rect 102086 711322 102322 711558
rect 102086 711002 102322 711238
rect 98386 709402 98622 709638
rect 98386 709082 98622 709318
rect 94686 707482 94922 707718
rect 94686 707162 94922 707398
rect 84086 697158 84322 697394
rect 84086 661158 84322 661394
rect 84086 625158 84322 625394
rect 84086 589158 84322 589394
rect 84086 553158 84322 553394
rect 84086 517158 84322 517394
rect 84086 481158 84322 481394
rect 84086 445158 84322 445394
rect 90986 705562 91222 705798
rect 90986 705242 91222 705478
rect 90986 668058 91222 668294
rect 90986 632058 91222 632294
rect 90986 596058 91222 596294
rect 90986 560058 91222 560294
rect 90986 524058 91222 524294
rect 90986 488058 91222 488294
rect 90986 452058 91222 452294
rect 94686 671758 94922 671994
rect 94686 635758 94922 635994
rect 94686 599758 94922 599994
rect 94686 563758 94922 563994
rect 94686 527758 94922 527994
rect 94686 491758 94922 491994
rect 94686 455758 94922 455994
rect 98386 675458 98622 675694
rect 98386 639458 98622 639694
rect 98386 603458 98622 603694
rect 98386 567458 98622 567694
rect 98386 531458 98622 531694
rect 98386 495458 98622 495694
rect 98386 459458 98622 459694
rect 120086 710362 120322 710598
rect 120086 710042 120322 710278
rect 116386 708442 116622 708678
rect 116386 708122 116622 708358
rect 112686 706522 112922 706758
rect 112686 706202 112922 706438
rect 102086 679158 102322 679394
rect 102086 643158 102322 643394
rect 102086 607158 102322 607394
rect 102086 571158 102322 571394
rect 102086 535158 102322 535394
rect 102086 499158 102322 499394
rect 102086 463158 102322 463394
rect 102086 427158 102322 427394
rect 108986 704602 109222 704838
rect 108986 704282 109222 704518
rect 108986 686058 109222 686294
rect 108986 650058 109222 650294
rect 108986 614058 109222 614294
rect 108986 578058 109222 578294
rect 108986 542058 109222 542294
rect 108986 506058 109222 506294
rect 108986 470058 109222 470294
rect 108986 434058 109222 434294
rect 112686 689758 112922 689994
rect 112686 653758 112922 653994
rect 112686 617758 112922 617994
rect 112686 581758 112922 581994
rect 112686 545758 112922 545994
rect 112686 509758 112922 509994
rect 112686 473758 112922 473994
rect 112686 437758 112922 437994
rect 116386 693458 116622 693694
rect 116386 657458 116622 657694
rect 116386 621458 116622 621694
rect 116386 585458 116622 585694
rect 116386 549458 116622 549694
rect 116386 513458 116622 513694
rect 116386 477458 116622 477694
rect 116386 441458 116622 441694
rect 138086 711322 138322 711558
rect 138086 711002 138322 711238
rect 134386 709402 134622 709638
rect 134386 709082 134622 709318
rect 130686 707482 130922 707718
rect 130686 707162 130922 707398
rect 120086 697158 120322 697394
rect 120086 661158 120322 661394
rect 120086 625158 120322 625394
rect 120086 589158 120322 589394
rect 120086 553158 120322 553394
rect 120086 517158 120322 517394
rect 120086 481158 120322 481394
rect 120086 445158 120322 445394
rect 126986 705562 127222 705798
rect 126986 705242 127222 705478
rect 126986 668058 127222 668294
rect 126986 632058 127222 632294
rect 126986 596058 127222 596294
rect 126986 560058 127222 560294
rect 126986 524058 127222 524294
rect 126986 488058 127222 488294
rect 126986 452058 127222 452294
rect 130686 671758 130922 671994
rect 130686 635758 130922 635994
rect 130686 599758 130922 599994
rect 130686 563758 130922 563994
rect 130686 527758 130922 527994
rect 130686 491758 130922 491994
rect 130686 455758 130922 455994
rect 134386 675458 134622 675694
rect 134386 639458 134622 639694
rect 134386 603458 134622 603694
rect 134386 567458 134622 567694
rect 134386 531458 134622 531694
rect 134386 495458 134622 495694
rect 134386 459458 134622 459694
rect 156086 710362 156322 710598
rect 156086 710042 156322 710278
rect 152386 708442 152622 708678
rect 152386 708122 152622 708358
rect 148686 706522 148922 706758
rect 148686 706202 148922 706438
rect 138086 679158 138322 679394
rect 138086 643158 138322 643394
rect 138086 607158 138322 607394
rect 138086 571158 138322 571394
rect 138086 535158 138322 535394
rect 138086 499158 138322 499394
rect 138086 463158 138322 463394
rect 138086 427158 138322 427394
rect 144986 704602 145222 704838
rect 144986 704282 145222 704518
rect 144986 686058 145222 686294
rect 144986 650058 145222 650294
rect 144986 614058 145222 614294
rect 144986 578058 145222 578294
rect 144986 542058 145222 542294
rect 144986 506058 145222 506294
rect 144986 470058 145222 470294
rect 144986 434058 145222 434294
rect 148686 689758 148922 689994
rect 148686 653758 148922 653994
rect 148686 617758 148922 617994
rect 148686 581758 148922 581994
rect 148686 545758 148922 545994
rect 148686 509758 148922 509994
rect 148686 473758 148922 473994
rect 148686 437758 148922 437994
rect 152386 693458 152622 693694
rect 152386 657458 152622 657694
rect 152386 621458 152622 621694
rect 152386 585458 152622 585694
rect 152386 549458 152622 549694
rect 152386 513458 152622 513694
rect 152386 477458 152622 477694
rect 152386 441458 152622 441694
rect 174086 711322 174322 711558
rect 174086 711002 174322 711238
rect 170386 709402 170622 709638
rect 170386 709082 170622 709318
rect 166686 707482 166922 707718
rect 166686 707162 166922 707398
rect 156086 697158 156322 697394
rect 156086 661158 156322 661394
rect 156086 625158 156322 625394
rect 156086 589158 156322 589394
rect 156086 553158 156322 553394
rect 156086 517158 156322 517394
rect 156086 481158 156322 481394
rect 156086 445158 156322 445394
rect 162986 705562 163222 705798
rect 162986 705242 163222 705478
rect 162986 668058 163222 668294
rect 162986 632058 163222 632294
rect 162986 596058 163222 596294
rect 162986 560058 163222 560294
rect 162986 524058 163222 524294
rect 162986 488058 163222 488294
rect 162986 452058 163222 452294
rect 166686 671758 166922 671994
rect 166686 635758 166922 635994
rect 166686 599758 166922 599994
rect 166686 563758 166922 563994
rect 166686 527758 166922 527994
rect 166686 491758 166922 491994
rect 166686 455758 166922 455994
rect 170386 675458 170622 675694
rect 170386 639458 170622 639694
rect 170386 603458 170622 603694
rect 170386 567458 170622 567694
rect 170386 531458 170622 531694
rect 170386 495458 170622 495694
rect 170386 459458 170622 459694
rect 192086 710362 192322 710598
rect 192086 710042 192322 710278
rect 188386 708442 188622 708678
rect 188386 708122 188622 708358
rect 184686 706522 184922 706758
rect 184686 706202 184922 706438
rect 174086 679158 174322 679394
rect 174086 643158 174322 643394
rect 174086 607158 174322 607394
rect 174086 571158 174322 571394
rect 174086 535158 174322 535394
rect 174086 499158 174322 499394
rect 174086 463158 174322 463394
rect 174086 427158 174322 427394
rect 180986 704602 181222 704838
rect 180986 704282 181222 704518
rect 180986 686058 181222 686294
rect 180986 650058 181222 650294
rect 180986 614058 181222 614294
rect 180986 578058 181222 578294
rect 180986 542058 181222 542294
rect 180986 506058 181222 506294
rect 180986 470058 181222 470294
rect 180986 434058 181222 434294
rect 40328 416058 40564 416294
rect 176056 416058 176292 416294
rect 36986 398058 37222 398294
rect 41008 398058 41244 398294
rect 175376 398058 175612 398294
rect 180986 398058 181222 398294
rect 40328 380058 40564 380294
rect 176056 380058 176292 380294
rect 36986 362058 37222 362294
rect 41008 362058 41244 362294
rect 175376 362058 175612 362294
rect 180986 362058 181222 362294
rect 40328 344058 40564 344294
rect 176056 344058 176292 344294
rect 36986 326058 37222 326294
rect 36986 290058 37222 290294
rect 36986 254058 37222 254294
rect 40686 329758 40922 329994
rect 40686 293758 40922 293994
rect 40686 257758 40922 257994
rect 44386 333458 44622 333694
rect 44386 297458 44622 297694
rect 44386 261458 44622 261694
rect 36986 218058 37222 218294
rect 36986 182058 37222 182294
rect 36986 146058 37222 146294
rect 36986 110058 37222 110294
rect 36986 74058 37222 74294
rect 44250 218058 44486 218294
rect 44250 182058 44486 182294
rect 44250 146058 44486 146294
rect 44250 110058 44486 110294
rect 44250 74058 44486 74294
rect 48086 337158 48322 337394
rect 48086 301158 48322 301394
rect 48086 265158 48322 265394
rect 54986 308058 55222 308294
rect 54986 272058 55222 272294
rect 58686 311758 58922 311994
rect 58686 275758 58922 275994
rect 62386 315458 62622 315694
rect 62386 279458 62622 279694
rect 66086 319158 66322 319394
rect 66086 283158 66322 283394
rect 66086 247158 66322 247394
rect 72986 326058 73222 326294
rect 72986 290058 73222 290294
rect 72986 254058 73222 254294
rect 76686 329758 76922 329994
rect 76686 293758 76922 293994
rect 76686 257758 76922 257994
rect 84086 337158 84322 337394
rect 80386 333458 80622 333694
rect 80386 297458 80622 297694
rect 80386 261458 80622 261694
rect 84086 301158 84322 301394
rect 84086 265158 84322 265394
rect 90986 308058 91222 308294
rect 90986 272058 91222 272294
rect 94686 311758 94922 311994
rect 94686 275758 94922 275994
rect 98386 315458 98622 315694
rect 98386 279458 98622 279694
rect 102086 319158 102322 319394
rect 102086 283158 102322 283394
rect 102086 247158 102322 247394
rect 108986 326058 109222 326294
rect 108986 290058 109222 290294
rect 108986 254058 109222 254294
rect 112686 329758 112922 329994
rect 112686 293758 112922 293994
rect 112686 257758 112922 257994
rect 116386 333458 116622 333694
rect 116386 297458 116622 297694
rect 116386 261458 116622 261694
rect 120086 337158 120322 337394
rect 120086 301158 120322 301394
rect 120086 265158 120322 265394
rect 126986 308058 127222 308294
rect 126986 272058 127222 272294
rect 130686 311758 130922 311994
rect 130686 275758 130922 275994
rect 134386 315458 134622 315694
rect 134386 279458 134622 279694
rect 138086 319158 138322 319394
rect 138086 283158 138322 283394
rect 138086 247158 138322 247394
rect 144986 326058 145222 326294
rect 144986 290058 145222 290294
rect 144986 254058 145222 254294
rect 148686 329758 148922 329994
rect 148686 293758 148922 293994
rect 148686 257758 148922 257994
rect 152386 333458 152622 333694
rect 152386 297458 152622 297694
rect 152386 261458 152622 261694
rect 156086 337158 156322 337394
rect 156086 301158 156322 301394
rect 156086 265158 156322 265394
rect 162986 308058 163222 308294
rect 162986 272058 163222 272294
rect 166686 311758 166922 311994
rect 166686 275758 166922 275994
rect 170386 315458 170622 315694
rect 170386 279458 170622 279694
rect 174086 319158 174322 319394
rect 174086 283158 174322 283394
rect 174086 247158 174322 247394
rect 180986 326058 181222 326294
rect 180986 290058 181222 290294
rect 180986 254058 181222 254294
rect 184686 689758 184922 689994
rect 184686 653758 184922 653994
rect 184686 617758 184922 617994
rect 184686 581758 184922 581994
rect 184686 545758 184922 545994
rect 184686 509758 184922 509994
rect 184686 473758 184922 473994
rect 184686 437758 184922 437994
rect 184686 401758 184922 401994
rect 184686 365758 184922 365994
rect 184686 329758 184922 329994
rect 184686 293758 184922 293994
rect 184686 257758 184922 257994
rect 188386 693458 188622 693694
rect 188386 657458 188622 657694
rect 188386 621458 188622 621694
rect 188386 585458 188622 585694
rect 188386 549458 188622 549694
rect 188386 513458 188622 513694
rect 188386 477458 188622 477694
rect 188386 441458 188622 441694
rect 188386 405458 188622 405694
rect 188386 369458 188622 369694
rect 188386 333458 188622 333694
rect 188386 297458 188622 297694
rect 188386 261458 188622 261694
rect 210086 711322 210322 711558
rect 210086 711002 210322 711238
rect 206386 709402 206622 709638
rect 206386 709082 206622 709318
rect 202686 707482 202922 707718
rect 202686 707162 202922 707398
rect 192086 697158 192322 697394
rect 192086 661158 192322 661394
rect 192086 625158 192322 625394
rect 192086 589158 192322 589394
rect 192086 553158 192322 553394
rect 192086 517158 192322 517394
rect 192086 481158 192322 481394
rect 192086 445158 192322 445394
rect 192086 409158 192322 409394
rect 192086 373158 192322 373394
rect 192086 337158 192322 337394
rect 192086 301158 192322 301394
rect 192086 265158 192322 265394
rect 198986 705562 199222 705798
rect 198986 705242 199222 705478
rect 198986 668058 199222 668294
rect 198986 632058 199222 632294
rect 198986 596058 199222 596294
rect 198986 560058 199222 560294
rect 198986 524058 199222 524294
rect 198986 488058 199222 488294
rect 198986 452058 199222 452294
rect 198986 416058 199222 416294
rect 198986 380058 199222 380294
rect 198986 344058 199222 344294
rect 198986 308058 199222 308294
rect 198986 272058 199222 272294
rect 202686 671758 202922 671994
rect 202686 635758 202922 635994
rect 202686 599758 202922 599994
rect 202686 563758 202922 563994
rect 202686 527758 202922 527994
rect 202686 491758 202922 491994
rect 202686 455758 202922 455994
rect 202686 419758 202922 419994
rect 202686 383758 202922 383994
rect 202686 347758 202922 347994
rect 202686 311758 202922 311994
rect 202686 275758 202922 275994
rect 206386 675458 206622 675694
rect 206386 639458 206622 639694
rect 206386 603458 206622 603694
rect 206386 567458 206622 567694
rect 206386 531458 206622 531694
rect 206386 495458 206622 495694
rect 206386 459458 206622 459694
rect 206386 423458 206622 423694
rect 206386 387458 206622 387694
rect 206386 351458 206622 351694
rect 206386 315458 206622 315694
rect 206386 279458 206622 279694
rect 228086 710362 228322 710598
rect 228086 710042 228322 710278
rect 224386 708442 224622 708678
rect 224386 708122 224622 708358
rect 220686 706522 220922 706758
rect 220686 706202 220922 706438
rect 210086 679158 210322 679394
rect 210086 643158 210322 643394
rect 210086 607158 210322 607394
rect 210086 571158 210322 571394
rect 210086 535158 210322 535394
rect 210086 499158 210322 499394
rect 210086 463158 210322 463394
rect 210086 427158 210322 427394
rect 210086 391158 210322 391394
rect 210086 355158 210322 355394
rect 210086 319158 210322 319394
rect 210086 283158 210322 283394
rect 210086 247158 210322 247394
rect 216986 704602 217222 704838
rect 216986 704282 217222 704518
rect 216986 686058 217222 686294
rect 216986 650058 217222 650294
rect 216986 614058 217222 614294
rect 216986 578058 217222 578294
rect 216986 542058 217222 542294
rect 216986 506058 217222 506294
rect 216986 470058 217222 470294
rect 216986 434058 217222 434294
rect 216986 398058 217222 398294
rect 216986 362058 217222 362294
rect 216986 326058 217222 326294
rect 216986 290058 217222 290294
rect 216986 254058 217222 254294
rect 220686 689758 220922 689994
rect 220686 653758 220922 653994
rect 220686 617758 220922 617994
rect 220686 581758 220922 581994
rect 220686 545758 220922 545994
rect 220686 509758 220922 509994
rect 220686 473758 220922 473994
rect 220686 437758 220922 437994
rect 220686 401758 220922 401994
rect 220686 365758 220922 365994
rect 220686 329758 220922 329994
rect 220686 293758 220922 293994
rect 220686 257758 220922 257994
rect 224386 693458 224622 693694
rect 224386 657458 224622 657694
rect 224386 621458 224622 621694
rect 224386 585458 224622 585694
rect 224386 549458 224622 549694
rect 224386 513458 224622 513694
rect 224386 477458 224622 477694
rect 224386 441458 224622 441694
rect 224386 405458 224622 405694
rect 224386 369458 224622 369694
rect 224386 333458 224622 333694
rect 224386 297458 224622 297694
rect 224386 261458 224622 261694
rect 246086 711322 246322 711558
rect 246086 711002 246322 711238
rect 242386 709402 242622 709638
rect 242386 709082 242622 709318
rect 238686 707482 238922 707718
rect 238686 707162 238922 707398
rect 228086 697158 228322 697394
rect 228086 661158 228322 661394
rect 228086 625158 228322 625394
rect 228086 589158 228322 589394
rect 228086 553158 228322 553394
rect 228086 517158 228322 517394
rect 228086 481158 228322 481394
rect 228086 445158 228322 445394
rect 228086 409158 228322 409394
rect 228086 373158 228322 373394
rect 228086 337158 228322 337394
rect 228086 301158 228322 301394
rect 228086 265158 228322 265394
rect 234986 705562 235222 705798
rect 234986 705242 235222 705478
rect 234986 668058 235222 668294
rect 234986 632058 235222 632294
rect 234986 596058 235222 596294
rect 234986 560058 235222 560294
rect 234986 524058 235222 524294
rect 234986 488058 235222 488294
rect 234986 452058 235222 452294
rect 234986 416058 235222 416294
rect 234986 380058 235222 380294
rect 234986 344058 235222 344294
rect 238686 671758 238922 671994
rect 238686 635758 238922 635994
rect 238686 599758 238922 599994
rect 238686 563758 238922 563994
rect 238686 527758 238922 527994
rect 238686 491758 238922 491994
rect 238686 455758 238922 455994
rect 238686 419758 238922 419994
rect 238686 383758 238922 383994
rect 238686 347758 238922 347994
rect 234986 308058 235222 308294
rect 234986 272058 235222 272294
rect 59610 236058 59846 236294
rect 90330 236058 90566 236294
rect 121050 236058 121286 236294
rect 151770 236058 152006 236294
rect 182490 236058 182726 236294
rect 213210 236058 213446 236294
rect 74970 218058 75206 218294
rect 105690 218058 105926 218294
rect 136410 218058 136646 218294
rect 167130 218058 167366 218294
rect 197850 218058 198086 218294
rect 228570 218058 228806 218294
rect 59610 200058 59846 200294
rect 90330 200058 90566 200294
rect 121050 200058 121286 200294
rect 151770 200058 152006 200294
rect 182490 200058 182726 200294
rect 213210 200058 213446 200294
rect 74970 182058 75206 182294
rect 105690 182058 105926 182294
rect 136410 182058 136646 182294
rect 167130 182058 167366 182294
rect 197850 182058 198086 182294
rect 228570 182058 228806 182294
rect 59610 164058 59846 164294
rect 90330 164058 90566 164294
rect 121050 164058 121286 164294
rect 151770 164058 152006 164294
rect 182490 164058 182726 164294
rect 213210 164058 213446 164294
rect 74970 146058 75206 146294
rect 105690 146058 105926 146294
rect 136410 146058 136646 146294
rect 167130 146058 167366 146294
rect 197850 146058 198086 146294
rect 228570 146058 228806 146294
rect 59610 128058 59846 128294
rect 90330 128058 90566 128294
rect 121050 128058 121286 128294
rect 151770 128058 152006 128294
rect 182490 128058 182726 128294
rect 213210 128058 213446 128294
rect 74970 110058 75206 110294
rect 105690 110058 105926 110294
rect 136410 110058 136646 110294
rect 167130 110058 167366 110294
rect 197850 110058 198086 110294
rect 228570 110058 228806 110294
rect 59610 92058 59846 92294
rect 90330 92058 90566 92294
rect 121050 92058 121286 92294
rect 151770 92058 152006 92294
rect 182490 92058 182726 92294
rect 213210 92058 213446 92294
rect 74970 74058 75206 74294
rect 105690 74058 105926 74294
rect 136410 74058 136646 74294
rect 167130 74058 167366 74294
rect 197850 74058 198086 74294
rect 228570 74058 228806 74294
rect 59610 56058 59846 56294
rect 90330 56058 90566 56294
rect 121050 56058 121286 56294
rect 151770 56058 152006 56294
rect 182490 56058 182726 56294
rect 213210 56058 213446 56294
rect 36986 38058 37222 38294
rect 36986 2058 37222 2294
rect 36986 -582 37222 -346
rect 36986 -902 37222 -666
rect 238686 311758 238922 311994
rect 238686 275758 238922 275994
rect 242386 675458 242622 675694
rect 242386 639458 242622 639694
rect 242386 603458 242622 603694
rect 242386 567458 242622 567694
rect 242386 531458 242622 531694
rect 242386 495458 242622 495694
rect 242386 459458 242622 459694
rect 242386 423458 242622 423694
rect 242386 387458 242622 387694
rect 242386 351458 242622 351694
rect 242386 315458 242622 315694
rect 242386 279458 242622 279694
rect 242386 243458 242622 243694
rect 242386 207458 242622 207694
rect 242386 171458 242622 171694
rect 242386 135458 242622 135694
rect 242386 99458 242622 99694
rect 242386 63458 242622 63694
rect 44386 9458 44622 9694
rect 40686 5758 40922 5994
rect 40686 -2502 40922 -2266
rect 40686 -2822 40922 -2586
rect 44386 -4422 44622 -4186
rect 44386 -4742 44622 -4506
rect 48086 13158 48322 13394
rect 30086 -7302 30322 -7066
rect 30086 -7622 30322 -7386
rect 54986 20058 55222 20294
rect 54986 -1542 55222 -1306
rect 54986 -1862 55222 -1626
rect 58686 23758 58922 23994
rect 58686 -3462 58922 -3226
rect 58686 -3782 58922 -3546
rect 62386 27458 62622 27694
rect 62386 -5382 62622 -5146
rect 62386 -5702 62622 -5466
rect 66086 31158 66322 31394
rect 48086 -6342 48322 -6106
rect 48086 -6662 48322 -6426
rect 72986 2058 73222 2294
rect 72986 -582 73222 -346
rect 72986 -902 73222 -666
rect 76686 5758 76922 5994
rect 76686 -2502 76922 -2266
rect 76686 -2822 76922 -2586
rect 80386 9458 80622 9694
rect 80386 -4422 80622 -4186
rect 80386 -4742 80622 -4506
rect 84086 13158 84322 13394
rect 66086 -7302 66322 -7066
rect 66086 -7622 66322 -7386
rect 90986 20058 91222 20294
rect 90986 -1542 91222 -1306
rect 90986 -1862 91222 -1626
rect 94686 23758 94922 23994
rect 94686 -3462 94922 -3226
rect 94686 -3782 94922 -3546
rect 98386 27458 98622 27694
rect 98386 -5382 98622 -5146
rect 98386 -5702 98622 -5466
rect 102086 31158 102322 31394
rect 84086 -6342 84322 -6106
rect 84086 -6662 84322 -6426
rect 108986 2058 109222 2294
rect 108986 -582 109222 -346
rect 108986 -902 109222 -666
rect 112686 5758 112922 5994
rect 112686 -2502 112922 -2266
rect 112686 -2822 112922 -2586
rect 116386 9458 116622 9694
rect 116386 -4422 116622 -4186
rect 116386 -4742 116622 -4506
rect 120086 13158 120322 13394
rect 102086 -7302 102322 -7066
rect 102086 -7622 102322 -7386
rect 126986 20058 127222 20294
rect 126986 -1542 127222 -1306
rect 126986 -1862 127222 -1626
rect 130686 23758 130922 23994
rect 130686 -3462 130922 -3226
rect 130686 -3782 130922 -3546
rect 134386 27458 134622 27694
rect 134386 -5382 134622 -5146
rect 134386 -5702 134622 -5466
rect 138086 31158 138322 31394
rect 120086 -6342 120322 -6106
rect 120086 -6662 120322 -6426
rect 144986 2058 145222 2294
rect 144986 -582 145222 -346
rect 144986 -902 145222 -666
rect 148686 5758 148922 5994
rect 148686 -2502 148922 -2266
rect 148686 -2822 148922 -2586
rect 152386 9458 152622 9694
rect 152386 -4422 152622 -4186
rect 152386 -4742 152622 -4506
rect 156086 13158 156322 13394
rect 138086 -7302 138322 -7066
rect 138086 -7622 138322 -7386
rect 162986 20058 163222 20294
rect 162986 -1542 163222 -1306
rect 162986 -1862 163222 -1626
rect 166686 23758 166922 23994
rect 166686 -3462 166922 -3226
rect 166686 -3782 166922 -3546
rect 170386 27458 170622 27694
rect 170386 -5382 170622 -5146
rect 170386 -5702 170622 -5466
rect 174086 31158 174322 31394
rect 156086 -6342 156322 -6106
rect 156086 -6662 156322 -6426
rect 180986 2058 181222 2294
rect 180986 -582 181222 -346
rect 180986 -902 181222 -666
rect 184686 5758 184922 5994
rect 184686 -2502 184922 -2266
rect 184686 -2822 184922 -2586
rect 188386 9458 188622 9694
rect 188386 -4422 188622 -4186
rect 188386 -4742 188622 -4506
rect 192086 13158 192322 13394
rect 174086 -7302 174322 -7066
rect 174086 -7622 174322 -7386
rect 198986 20058 199222 20294
rect 198986 -1542 199222 -1306
rect 198986 -1862 199222 -1626
rect 202686 23758 202922 23994
rect 202686 -3462 202922 -3226
rect 202686 -3782 202922 -3546
rect 206386 27458 206622 27694
rect 206386 -5382 206622 -5146
rect 206386 -5702 206622 -5466
rect 210086 31158 210322 31394
rect 192086 -6342 192322 -6106
rect 192086 -6662 192322 -6426
rect 216986 2058 217222 2294
rect 216986 -582 217222 -346
rect 216986 -902 217222 -666
rect 220686 5758 220922 5994
rect 220686 -2502 220922 -2266
rect 220686 -2822 220922 -2586
rect 224386 9458 224622 9694
rect 224386 -4422 224622 -4186
rect 224386 -4742 224622 -4506
rect 228086 13158 228322 13394
rect 210086 -7302 210322 -7066
rect 210086 -7622 210322 -7386
rect 234986 20058 235222 20294
rect 234986 -1542 235222 -1306
rect 234986 -1862 235222 -1626
rect 238686 23758 238922 23994
rect 238686 -3462 238922 -3226
rect 238686 -3782 238922 -3546
rect 242386 27458 242622 27694
rect 242386 -5382 242622 -5146
rect 242386 -5702 242622 -5466
rect 264086 710362 264322 710598
rect 264086 710042 264322 710278
rect 260386 708442 260622 708678
rect 260386 708122 260622 708358
rect 256686 706522 256922 706758
rect 256686 706202 256922 706438
rect 246086 679158 246322 679394
rect 246086 643158 246322 643394
rect 246086 607158 246322 607394
rect 246086 571158 246322 571394
rect 246086 535158 246322 535394
rect 246086 499158 246322 499394
rect 246086 463158 246322 463394
rect 246086 427158 246322 427394
rect 246086 391158 246322 391394
rect 246086 355158 246322 355394
rect 246086 319158 246322 319394
rect 246086 283158 246322 283394
rect 246086 247158 246322 247394
rect 246086 211158 246322 211394
rect 246086 175158 246322 175394
rect 246086 139158 246322 139394
rect 246086 103158 246322 103394
rect 246086 67158 246322 67394
rect 246086 31158 246322 31394
rect 228086 -6342 228322 -6106
rect 228086 -6662 228322 -6426
rect 252986 704602 253222 704838
rect 252986 704282 253222 704518
rect 252986 686058 253222 686294
rect 252986 650058 253222 650294
rect 252986 614058 253222 614294
rect 252986 578058 253222 578294
rect 252986 542058 253222 542294
rect 252986 506058 253222 506294
rect 252986 470058 253222 470294
rect 252986 434058 253222 434294
rect 252986 398058 253222 398294
rect 252986 362058 253222 362294
rect 252986 326058 253222 326294
rect 252986 290058 253222 290294
rect 252986 254058 253222 254294
rect 252986 218058 253222 218294
rect 252986 182058 253222 182294
rect 252986 146058 253222 146294
rect 252986 110058 253222 110294
rect 252986 74058 253222 74294
rect 252986 38058 253222 38294
rect 252986 2058 253222 2294
rect 252986 -582 253222 -346
rect 252986 -902 253222 -666
rect 256686 689758 256922 689994
rect 256686 653758 256922 653994
rect 256686 617758 256922 617994
rect 256686 581758 256922 581994
rect 256686 545758 256922 545994
rect 256686 509758 256922 509994
rect 256686 473758 256922 473994
rect 256686 437758 256922 437994
rect 256686 401758 256922 401994
rect 256686 365758 256922 365994
rect 256686 329758 256922 329994
rect 256686 293758 256922 293994
rect 256686 257758 256922 257994
rect 256686 221758 256922 221994
rect 256686 185758 256922 185994
rect 256686 149758 256922 149994
rect 256686 113758 256922 113994
rect 256686 77758 256922 77994
rect 256686 41758 256922 41994
rect 256686 5758 256922 5994
rect 256686 -2502 256922 -2266
rect 256686 -2822 256922 -2586
rect 260386 693458 260622 693694
rect 260386 657458 260622 657694
rect 260386 621458 260622 621694
rect 260386 585458 260622 585694
rect 260386 549458 260622 549694
rect 260386 513458 260622 513694
rect 260386 477458 260622 477694
rect 260386 441458 260622 441694
rect 260386 405458 260622 405694
rect 260386 369458 260622 369694
rect 260386 333458 260622 333694
rect 260386 297458 260622 297694
rect 260386 261458 260622 261694
rect 260386 225458 260622 225694
rect 260386 189458 260622 189694
rect 260386 153458 260622 153694
rect 260386 117458 260622 117694
rect 260386 81458 260622 81694
rect 260386 45458 260622 45694
rect 260386 9458 260622 9694
rect 260386 -4422 260622 -4186
rect 260386 -4742 260622 -4506
rect 282086 711322 282322 711558
rect 282086 711002 282322 711238
rect 278386 709402 278622 709638
rect 278386 709082 278622 709318
rect 274686 707482 274922 707718
rect 274686 707162 274922 707398
rect 264086 697158 264322 697394
rect 264086 661158 264322 661394
rect 264086 625158 264322 625394
rect 264086 589158 264322 589394
rect 264086 553158 264322 553394
rect 264086 517158 264322 517394
rect 264086 481158 264322 481394
rect 264086 445158 264322 445394
rect 264086 409158 264322 409394
rect 264086 373158 264322 373394
rect 264086 337158 264322 337394
rect 264086 301158 264322 301394
rect 264086 265158 264322 265394
rect 264086 229158 264322 229394
rect 264086 193158 264322 193394
rect 264086 157158 264322 157394
rect 264086 121158 264322 121394
rect 264086 85158 264322 85394
rect 264086 49158 264322 49394
rect 264086 13158 264322 13394
rect 246086 -7302 246322 -7066
rect 246086 -7622 246322 -7386
rect 270986 705562 271222 705798
rect 270986 705242 271222 705478
rect 270986 668058 271222 668294
rect 270986 632058 271222 632294
rect 270986 596058 271222 596294
rect 270986 560058 271222 560294
rect 270986 524058 271222 524294
rect 270986 488058 271222 488294
rect 270986 452058 271222 452294
rect 270986 416058 271222 416294
rect 270986 380058 271222 380294
rect 270986 344058 271222 344294
rect 270986 308058 271222 308294
rect 270986 272058 271222 272294
rect 270986 236058 271222 236294
rect 270986 200058 271222 200294
rect 270986 164058 271222 164294
rect 270986 128058 271222 128294
rect 270986 92058 271222 92294
rect 270986 56058 271222 56294
rect 270986 20058 271222 20294
rect 270986 -1542 271222 -1306
rect 270986 -1862 271222 -1626
rect 274686 671758 274922 671994
rect 274686 635758 274922 635994
rect 274686 599758 274922 599994
rect 274686 563758 274922 563994
rect 274686 527758 274922 527994
rect 274686 491758 274922 491994
rect 274686 455758 274922 455994
rect 274686 419758 274922 419994
rect 274686 383758 274922 383994
rect 274686 347758 274922 347994
rect 274686 311758 274922 311994
rect 274686 275758 274922 275994
rect 274686 239758 274922 239994
rect 274686 203758 274922 203994
rect 274686 167758 274922 167994
rect 274686 131758 274922 131994
rect 274686 95758 274922 95994
rect 274686 59758 274922 59994
rect 274686 23758 274922 23994
rect 274686 -3462 274922 -3226
rect 274686 -3782 274922 -3546
rect 278386 675458 278622 675694
rect 278386 639458 278622 639694
rect 278386 603458 278622 603694
rect 278386 567458 278622 567694
rect 278386 531458 278622 531694
rect 278386 495458 278622 495694
rect 278386 459458 278622 459694
rect 278386 423458 278622 423694
rect 278386 387458 278622 387694
rect 278386 351458 278622 351694
rect 278386 315458 278622 315694
rect 278386 279458 278622 279694
rect 278386 243458 278622 243694
rect 278386 207458 278622 207694
rect 278386 171458 278622 171694
rect 278386 135458 278622 135694
rect 278386 99458 278622 99694
rect 278386 63458 278622 63694
rect 278386 27458 278622 27694
rect 278386 -5382 278622 -5146
rect 278386 -5702 278622 -5466
rect 300086 710362 300322 710598
rect 300086 710042 300322 710278
rect 296386 708442 296622 708678
rect 296386 708122 296622 708358
rect 292686 706522 292922 706758
rect 292686 706202 292922 706438
rect 282086 679158 282322 679394
rect 282086 643158 282322 643394
rect 282086 607158 282322 607394
rect 282086 571158 282322 571394
rect 282086 535158 282322 535394
rect 282086 499158 282322 499394
rect 282086 463158 282322 463394
rect 282086 427158 282322 427394
rect 282086 391158 282322 391394
rect 282086 355158 282322 355394
rect 282086 319158 282322 319394
rect 282086 283158 282322 283394
rect 282086 247158 282322 247394
rect 282086 211158 282322 211394
rect 282086 175158 282322 175394
rect 282086 139158 282322 139394
rect 282086 103158 282322 103394
rect 282086 67158 282322 67394
rect 282086 31158 282322 31394
rect 264086 -6342 264322 -6106
rect 264086 -6662 264322 -6426
rect 288986 704602 289222 704838
rect 288986 704282 289222 704518
rect 288986 686058 289222 686294
rect 288986 650058 289222 650294
rect 288986 614058 289222 614294
rect 288986 578058 289222 578294
rect 288986 542058 289222 542294
rect 288986 506058 289222 506294
rect 288986 470058 289222 470294
rect 288986 434058 289222 434294
rect 288986 398058 289222 398294
rect 288986 362058 289222 362294
rect 288986 326058 289222 326294
rect 288986 290058 289222 290294
rect 288986 254058 289222 254294
rect 288986 218058 289222 218294
rect 288986 182058 289222 182294
rect 288986 146058 289222 146294
rect 288986 110058 289222 110294
rect 288986 74058 289222 74294
rect 288986 38058 289222 38294
rect 288986 2058 289222 2294
rect 288986 -582 289222 -346
rect 288986 -902 289222 -666
rect 292686 689758 292922 689994
rect 292686 653758 292922 653994
rect 292686 617758 292922 617994
rect 292686 581758 292922 581994
rect 292686 545758 292922 545994
rect 292686 509758 292922 509994
rect 292686 473758 292922 473994
rect 292686 437758 292922 437994
rect 292686 401758 292922 401994
rect 292686 365758 292922 365994
rect 292686 329758 292922 329994
rect 292686 293758 292922 293994
rect 292686 257758 292922 257994
rect 292686 221758 292922 221994
rect 292686 185758 292922 185994
rect 292686 149758 292922 149994
rect 292686 113758 292922 113994
rect 292686 77758 292922 77994
rect 292686 41758 292922 41994
rect 292686 5758 292922 5994
rect 292686 -2502 292922 -2266
rect 292686 -2822 292922 -2586
rect 296386 693458 296622 693694
rect 296386 657458 296622 657694
rect 296386 621458 296622 621694
rect 296386 585458 296622 585694
rect 296386 549458 296622 549694
rect 296386 513458 296622 513694
rect 296386 477458 296622 477694
rect 296386 441458 296622 441694
rect 296386 405458 296622 405694
rect 296386 369458 296622 369694
rect 296386 333458 296622 333694
rect 296386 297458 296622 297694
rect 296386 261458 296622 261694
rect 296386 225458 296622 225694
rect 296386 189458 296622 189694
rect 296386 153458 296622 153694
rect 296386 117458 296622 117694
rect 296386 81458 296622 81694
rect 296386 45458 296622 45694
rect 296386 9458 296622 9694
rect 296386 -4422 296622 -4186
rect 296386 -4742 296622 -4506
rect 318086 711322 318322 711558
rect 318086 711002 318322 711238
rect 314386 709402 314622 709638
rect 314386 709082 314622 709318
rect 310686 707482 310922 707718
rect 310686 707162 310922 707398
rect 300086 697158 300322 697394
rect 300086 661158 300322 661394
rect 300086 625158 300322 625394
rect 300086 589158 300322 589394
rect 300086 553158 300322 553394
rect 300086 517158 300322 517394
rect 300086 481158 300322 481394
rect 300086 445158 300322 445394
rect 300086 409158 300322 409394
rect 300086 373158 300322 373394
rect 300086 337158 300322 337394
rect 300086 301158 300322 301394
rect 300086 265158 300322 265394
rect 300086 229158 300322 229394
rect 300086 193158 300322 193394
rect 300086 157158 300322 157394
rect 300086 121158 300322 121394
rect 300086 85158 300322 85394
rect 300086 49158 300322 49394
rect 300086 13158 300322 13394
rect 282086 -7302 282322 -7066
rect 282086 -7622 282322 -7386
rect 306986 705562 307222 705798
rect 306986 705242 307222 705478
rect 306986 668058 307222 668294
rect 306986 632058 307222 632294
rect 306986 596058 307222 596294
rect 306986 560058 307222 560294
rect 306986 524058 307222 524294
rect 306986 488058 307222 488294
rect 306986 452058 307222 452294
rect 306986 416058 307222 416294
rect 306986 380058 307222 380294
rect 306986 344058 307222 344294
rect 306986 308058 307222 308294
rect 306986 272058 307222 272294
rect 306986 236058 307222 236294
rect 306986 200058 307222 200294
rect 306986 164058 307222 164294
rect 306986 128058 307222 128294
rect 306986 92058 307222 92294
rect 306986 56058 307222 56294
rect 306986 20058 307222 20294
rect 306986 -1542 307222 -1306
rect 306986 -1862 307222 -1626
rect 310686 671758 310922 671994
rect 310686 635758 310922 635994
rect 310686 599758 310922 599994
rect 310686 563758 310922 563994
rect 310686 527758 310922 527994
rect 310686 491758 310922 491994
rect 310686 455758 310922 455994
rect 310686 419758 310922 419994
rect 310686 383758 310922 383994
rect 310686 347758 310922 347994
rect 310686 311758 310922 311994
rect 310686 275758 310922 275994
rect 310686 239758 310922 239994
rect 310686 203758 310922 203994
rect 310686 167758 310922 167994
rect 310686 131758 310922 131994
rect 310686 95758 310922 95994
rect 310686 59758 310922 59994
rect 310686 23758 310922 23994
rect 310686 -3462 310922 -3226
rect 310686 -3782 310922 -3546
rect 314386 675458 314622 675694
rect 314386 639458 314622 639694
rect 314386 603458 314622 603694
rect 314386 567458 314622 567694
rect 314386 531458 314622 531694
rect 314386 495458 314622 495694
rect 314386 459458 314622 459694
rect 314386 423458 314622 423694
rect 314386 387458 314622 387694
rect 314386 351458 314622 351694
rect 314386 315458 314622 315694
rect 314386 279458 314622 279694
rect 314386 243458 314622 243694
rect 314386 207458 314622 207694
rect 314386 171458 314622 171694
rect 314386 135458 314622 135694
rect 314386 99458 314622 99694
rect 314386 63458 314622 63694
rect 314386 27458 314622 27694
rect 314386 -5382 314622 -5146
rect 314386 -5702 314622 -5466
rect 336086 710362 336322 710598
rect 336086 710042 336322 710278
rect 332386 708442 332622 708678
rect 332386 708122 332622 708358
rect 328686 706522 328922 706758
rect 328686 706202 328922 706438
rect 318086 679158 318322 679394
rect 318086 643158 318322 643394
rect 318086 607158 318322 607394
rect 318086 571158 318322 571394
rect 318086 535158 318322 535394
rect 318086 499158 318322 499394
rect 318086 463158 318322 463394
rect 318086 427158 318322 427394
rect 318086 391158 318322 391394
rect 318086 355158 318322 355394
rect 318086 319158 318322 319394
rect 318086 283158 318322 283394
rect 318086 247158 318322 247394
rect 318086 211158 318322 211394
rect 318086 175158 318322 175394
rect 318086 139158 318322 139394
rect 318086 103158 318322 103394
rect 318086 67158 318322 67394
rect 318086 31158 318322 31394
rect 300086 -6342 300322 -6106
rect 300086 -6662 300322 -6426
rect 324986 704602 325222 704838
rect 324986 704282 325222 704518
rect 324986 686058 325222 686294
rect 324986 650058 325222 650294
rect 324986 614058 325222 614294
rect 324986 578058 325222 578294
rect 324986 542058 325222 542294
rect 324986 506058 325222 506294
rect 324986 470058 325222 470294
rect 324986 434058 325222 434294
rect 324986 398058 325222 398294
rect 324986 362058 325222 362294
rect 324986 326058 325222 326294
rect 324986 290058 325222 290294
rect 324986 254058 325222 254294
rect 324986 218058 325222 218294
rect 324986 182058 325222 182294
rect 324986 146058 325222 146294
rect 324986 110058 325222 110294
rect 324986 74058 325222 74294
rect 324986 38058 325222 38294
rect 324986 2058 325222 2294
rect 324986 -582 325222 -346
rect 324986 -902 325222 -666
rect 328686 689758 328922 689994
rect 328686 653758 328922 653994
rect 328686 617758 328922 617994
rect 328686 581758 328922 581994
rect 328686 545758 328922 545994
rect 328686 509758 328922 509994
rect 328686 473758 328922 473994
rect 328686 437758 328922 437994
rect 328686 401758 328922 401994
rect 328686 365758 328922 365994
rect 328686 329758 328922 329994
rect 328686 293758 328922 293994
rect 328686 257758 328922 257994
rect 328686 221758 328922 221994
rect 328686 185758 328922 185994
rect 328686 149758 328922 149994
rect 328686 113758 328922 113994
rect 328686 77758 328922 77994
rect 328686 41758 328922 41994
rect 328686 5758 328922 5994
rect 328686 -2502 328922 -2266
rect 328686 -2822 328922 -2586
rect 332386 693458 332622 693694
rect 332386 657458 332622 657694
rect 332386 621458 332622 621694
rect 332386 585458 332622 585694
rect 332386 549458 332622 549694
rect 332386 513458 332622 513694
rect 332386 477458 332622 477694
rect 332386 441458 332622 441694
rect 332386 405458 332622 405694
rect 332386 369458 332622 369694
rect 332386 333458 332622 333694
rect 332386 297458 332622 297694
rect 332386 261458 332622 261694
rect 332386 225458 332622 225694
rect 332386 189458 332622 189694
rect 332386 153458 332622 153694
rect 332386 117458 332622 117694
rect 332386 81458 332622 81694
rect 332386 45458 332622 45694
rect 332386 9458 332622 9694
rect 332386 -4422 332622 -4186
rect 332386 -4742 332622 -4506
rect 354086 711322 354322 711558
rect 354086 711002 354322 711238
rect 350386 709402 350622 709638
rect 350386 709082 350622 709318
rect 346686 707482 346922 707718
rect 346686 707162 346922 707398
rect 336086 697158 336322 697394
rect 336086 661158 336322 661394
rect 336086 625158 336322 625394
rect 336086 589158 336322 589394
rect 336086 553158 336322 553394
rect 336086 517158 336322 517394
rect 336086 481158 336322 481394
rect 336086 445158 336322 445394
rect 342986 705562 343222 705798
rect 342986 705242 343222 705478
rect 342986 668058 343222 668294
rect 342986 632058 343222 632294
rect 342986 596058 343222 596294
rect 342986 560058 343222 560294
rect 342986 524058 343222 524294
rect 342986 488058 343222 488294
rect 342986 452058 343222 452294
rect 346686 671758 346922 671994
rect 346686 635758 346922 635994
rect 346686 599758 346922 599994
rect 346686 563758 346922 563994
rect 346686 527758 346922 527994
rect 346686 491758 346922 491994
rect 346686 455758 346922 455994
rect 350386 675458 350622 675694
rect 350386 639458 350622 639694
rect 350386 603458 350622 603694
rect 350386 567458 350622 567694
rect 350386 531458 350622 531694
rect 350386 495458 350622 495694
rect 350386 459458 350622 459694
rect 372086 710362 372322 710598
rect 372086 710042 372322 710278
rect 368386 708442 368622 708678
rect 368386 708122 368622 708358
rect 364686 706522 364922 706758
rect 364686 706202 364922 706438
rect 354086 679158 354322 679394
rect 354086 643158 354322 643394
rect 354086 607158 354322 607394
rect 354086 571158 354322 571394
rect 354086 535158 354322 535394
rect 354086 499158 354322 499394
rect 354086 463158 354322 463394
rect 354086 427158 354322 427394
rect 360986 704602 361222 704838
rect 360986 704282 361222 704518
rect 360986 686058 361222 686294
rect 360986 650058 361222 650294
rect 360986 614058 361222 614294
rect 360986 578058 361222 578294
rect 360986 542058 361222 542294
rect 360986 506058 361222 506294
rect 360986 470058 361222 470294
rect 360986 434058 361222 434294
rect 364686 689758 364922 689994
rect 364686 653758 364922 653994
rect 364686 617758 364922 617994
rect 364686 581758 364922 581994
rect 364686 545758 364922 545994
rect 364686 509758 364922 509994
rect 364686 473758 364922 473994
rect 364686 437758 364922 437994
rect 368386 693458 368622 693694
rect 368386 657458 368622 657694
rect 368386 621458 368622 621694
rect 368386 585458 368622 585694
rect 368386 549458 368622 549694
rect 368386 513458 368622 513694
rect 368386 477458 368622 477694
rect 368386 441458 368622 441694
rect 390086 711322 390322 711558
rect 390086 711002 390322 711238
rect 386386 709402 386622 709638
rect 386386 709082 386622 709318
rect 382686 707482 382922 707718
rect 382686 707162 382922 707398
rect 372086 697158 372322 697394
rect 372086 661158 372322 661394
rect 372086 625158 372322 625394
rect 372086 589158 372322 589394
rect 372086 553158 372322 553394
rect 372086 517158 372322 517394
rect 372086 481158 372322 481394
rect 372086 445158 372322 445394
rect 378986 705562 379222 705798
rect 378986 705242 379222 705478
rect 378986 668058 379222 668294
rect 378986 632058 379222 632294
rect 378986 596058 379222 596294
rect 378986 560058 379222 560294
rect 378986 524058 379222 524294
rect 378986 488058 379222 488294
rect 378986 452058 379222 452294
rect 382686 671758 382922 671994
rect 382686 635758 382922 635994
rect 382686 599758 382922 599994
rect 382686 563758 382922 563994
rect 382686 527758 382922 527994
rect 382686 491758 382922 491994
rect 382686 455758 382922 455994
rect 386386 675458 386622 675694
rect 386386 639458 386622 639694
rect 386386 603458 386622 603694
rect 386386 567458 386622 567694
rect 386386 531458 386622 531694
rect 386386 495458 386622 495694
rect 386386 459458 386622 459694
rect 408086 710362 408322 710598
rect 408086 710042 408322 710278
rect 404386 708442 404622 708678
rect 404386 708122 404622 708358
rect 400686 706522 400922 706758
rect 400686 706202 400922 706438
rect 390086 679158 390322 679394
rect 390086 643158 390322 643394
rect 390086 607158 390322 607394
rect 390086 571158 390322 571394
rect 390086 535158 390322 535394
rect 390086 499158 390322 499394
rect 390086 463158 390322 463394
rect 390086 427158 390322 427394
rect 396986 704602 397222 704838
rect 396986 704282 397222 704518
rect 396986 686058 397222 686294
rect 396986 650058 397222 650294
rect 396986 614058 397222 614294
rect 396986 578058 397222 578294
rect 396986 542058 397222 542294
rect 396986 506058 397222 506294
rect 396986 470058 397222 470294
rect 396986 434058 397222 434294
rect 400686 689758 400922 689994
rect 400686 653758 400922 653994
rect 400686 617758 400922 617994
rect 400686 581758 400922 581994
rect 400686 545758 400922 545994
rect 400686 509758 400922 509994
rect 400686 473758 400922 473994
rect 400686 437758 400922 437994
rect 404386 693458 404622 693694
rect 404386 657458 404622 657694
rect 404386 621458 404622 621694
rect 404386 585458 404622 585694
rect 404386 549458 404622 549694
rect 404386 513458 404622 513694
rect 404386 477458 404622 477694
rect 404386 441458 404622 441694
rect 426086 711322 426322 711558
rect 426086 711002 426322 711238
rect 422386 709402 422622 709638
rect 422386 709082 422622 709318
rect 418686 707482 418922 707718
rect 418686 707162 418922 707398
rect 408086 697158 408322 697394
rect 408086 661158 408322 661394
rect 408086 625158 408322 625394
rect 408086 589158 408322 589394
rect 408086 553158 408322 553394
rect 408086 517158 408322 517394
rect 408086 481158 408322 481394
rect 408086 445158 408322 445394
rect 414986 705562 415222 705798
rect 414986 705242 415222 705478
rect 414986 668058 415222 668294
rect 414986 632058 415222 632294
rect 414986 596058 415222 596294
rect 414986 560058 415222 560294
rect 414986 524058 415222 524294
rect 414986 488058 415222 488294
rect 414986 452058 415222 452294
rect 418686 671758 418922 671994
rect 418686 635758 418922 635994
rect 418686 599758 418922 599994
rect 418686 563758 418922 563994
rect 418686 527758 418922 527994
rect 418686 491758 418922 491994
rect 418686 455758 418922 455994
rect 422386 675458 422622 675694
rect 422386 639458 422622 639694
rect 422386 603458 422622 603694
rect 422386 567458 422622 567694
rect 422386 531458 422622 531694
rect 422386 495458 422622 495694
rect 422386 459458 422622 459694
rect 444086 710362 444322 710598
rect 444086 710042 444322 710278
rect 440386 708442 440622 708678
rect 440386 708122 440622 708358
rect 436686 706522 436922 706758
rect 436686 706202 436922 706438
rect 426086 679158 426322 679394
rect 426086 643158 426322 643394
rect 426086 607158 426322 607394
rect 426086 571158 426322 571394
rect 426086 535158 426322 535394
rect 426086 499158 426322 499394
rect 426086 463158 426322 463394
rect 426086 427158 426322 427394
rect 432986 704602 433222 704838
rect 432986 704282 433222 704518
rect 432986 686058 433222 686294
rect 432986 650058 433222 650294
rect 432986 614058 433222 614294
rect 432986 578058 433222 578294
rect 432986 542058 433222 542294
rect 432986 506058 433222 506294
rect 432986 470058 433222 470294
rect 432986 434058 433222 434294
rect 436686 689758 436922 689994
rect 436686 653758 436922 653994
rect 436686 617758 436922 617994
rect 436686 581758 436922 581994
rect 436686 545758 436922 545994
rect 436686 509758 436922 509994
rect 436686 473758 436922 473994
rect 436686 437758 436922 437994
rect 440386 693458 440622 693694
rect 440386 657458 440622 657694
rect 440386 621458 440622 621694
rect 440386 585458 440622 585694
rect 440386 549458 440622 549694
rect 440386 513458 440622 513694
rect 440386 477458 440622 477694
rect 440386 441458 440622 441694
rect 462086 711322 462322 711558
rect 462086 711002 462322 711238
rect 458386 709402 458622 709638
rect 458386 709082 458622 709318
rect 454686 707482 454922 707718
rect 454686 707162 454922 707398
rect 444086 697158 444322 697394
rect 444086 661158 444322 661394
rect 444086 625158 444322 625394
rect 444086 589158 444322 589394
rect 444086 553158 444322 553394
rect 444086 517158 444322 517394
rect 444086 481158 444322 481394
rect 444086 445158 444322 445394
rect 450986 705562 451222 705798
rect 450986 705242 451222 705478
rect 450986 668058 451222 668294
rect 450986 632058 451222 632294
rect 450986 596058 451222 596294
rect 450986 560058 451222 560294
rect 450986 524058 451222 524294
rect 450986 488058 451222 488294
rect 450986 452058 451222 452294
rect 454686 671758 454922 671994
rect 454686 635758 454922 635994
rect 454686 599758 454922 599994
rect 454686 563758 454922 563994
rect 454686 527758 454922 527994
rect 454686 491758 454922 491994
rect 454686 455758 454922 455994
rect 458386 675458 458622 675694
rect 458386 639458 458622 639694
rect 458386 603458 458622 603694
rect 458386 567458 458622 567694
rect 458386 531458 458622 531694
rect 458386 495458 458622 495694
rect 458386 459458 458622 459694
rect 480086 710362 480322 710598
rect 480086 710042 480322 710278
rect 476386 708442 476622 708678
rect 476386 708122 476622 708358
rect 472686 706522 472922 706758
rect 472686 706202 472922 706438
rect 462086 679158 462322 679394
rect 462086 643158 462322 643394
rect 462086 607158 462322 607394
rect 462086 571158 462322 571394
rect 462086 535158 462322 535394
rect 462086 499158 462322 499394
rect 462086 463158 462322 463394
rect 462086 427158 462322 427394
rect 468986 704602 469222 704838
rect 468986 704282 469222 704518
rect 468986 686058 469222 686294
rect 468986 650058 469222 650294
rect 468986 614058 469222 614294
rect 468986 578058 469222 578294
rect 468986 542058 469222 542294
rect 468986 506058 469222 506294
rect 468986 470058 469222 470294
rect 468986 434058 469222 434294
rect 472686 689758 472922 689994
rect 472686 653758 472922 653994
rect 472686 617758 472922 617994
rect 472686 581758 472922 581994
rect 472686 545758 472922 545994
rect 472686 509758 472922 509994
rect 472686 473758 472922 473994
rect 472686 437758 472922 437994
rect 476386 693458 476622 693694
rect 476386 657458 476622 657694
rect 476386 621458 476622 621694
rect 476386 585458 476622 585694
rect 476386 549458 476622 549694
rect 476386 513458 476622 513694
rect 476386 477458 476622 477694
rect 476386 441458 476622 441694
rect 498086 711322 498322 711558
rect 498086 711002 498322 711238
rect 494386 709402 494622 709638
rect 494386 709082 494622 709318
rect 490686 707482 490922 707718
rect 490686 707162 490922 707398
rect 480086 697158 480322 697394
rect 480086 661158 480322 661394
rect 480086 625158 480322 625394
rect 480086 589158 480322 589394
rect 480086 553158 480322 553394
rect 480086 517158 480322 517394
rect 480086 481158 480322 481394
rect 480086 445158 480322 445394
rect 340328 416058 340564 416294
rect 476056 416058 476292 416294
rect 336086 409158 336322 409394
rect 480086 409158 480322 409394
rect 341008 398058 341244 398294
rect 475376 398058 475612 398294
rect 340328 380058 340564 380294
rect 476056 380058 476292 380294
rect 336086 373158 336322 373394
rect 480086 373158 480322 373394
rect 341008 362058 341244 362294
rect 475376 362058 475612 362294
rect 340328 344058 340564 344294
rect 476056 344058 476292 344294
rect 336086 337158 336322 337394
rect 336086 301158 336322 301394
rect 336086 265158 336322 265394
rect 336086 229158 336322 229394
rect 336086 193158 336322 193394
rect 336086 157158 336322 157394
rect 336086 121158 336322 121394
rect 336086 85158 336322 85394
rect 336086 49158 336322 49394
rect 336086 13158 336322 13394
rect 318086 -7302 318322 -7066
rect 318086 -7622 318322 -7386
rect 342986 308058 343222 308294
rect 342986 272058 343222 272294
rect 342986 236058 343222 236294
rect 342986 200058 343222 200294
rect 342986 164058 343222 164294
rect 342986 128058 343222 128294
rect 342986 92058 343222 92294
rect 342986 56058 343222 56294
rect 342986 20058 343222 20294
rect 342986 -1542 343222 -1306
rect 342986 -1862 343222 -1626
rect 346686 311758 346922 311994
rect 346686 275758 346922 275994
rect 346686 239758 346922 239994
rect 346686 203758 346922 203994
rect 346686 167758 346922 167994
rect 346686 131758 346922 131994
rect 346686 95758 346922 95994
rect 346686 59758 346922 59994
rect 346686 23758 346922 23994
rect 346686 -3462 346922 -3226
rect 346686 -3782 346922 -3546
rect 350386 315458 350622 315694
rect 350386 279458 350622 279694
rect 350386 243458 350622 243694
rect 350386 207458 350622 207694
rect 350386 171458 350622 171694
rect 350386 135458 350622 135694
rect 350386 99458 350622 99694
rect 350386 63458 350622 63694
rect 350386 27458 350622 27694
rect 350386 -5382 350622 -5146
rect 350386 -5702 350622 -5466
rect 354086 319158 354322 319394
rect 354086 283158 354322 283394
rect 354086 247158 354322 247394
rect 354086 211158 354322 211394
rect 354086 175158 354322 175394
rect 354086 139158 354322 139394
rect 354086 103158 354322 103394
rect 354086 67158 354322 67394
rect 354086 31158 354322 31394
rect 336086 -6342 336322 -6106
rect 336086 -6662 336322 -6426
rect 360986 326058 361222 326294
rect 360986 290058 361222 290294
rect 360986 254058 361222 254294
rect 360986 218058 361222 218294
rect 360986 182058 361222 182294
rect 360986 146058 361222 146294
rect 360986 110058 361222 110294
rect 360986 74058 361222 74294
rect 360986 38058 361222 38294
rect 360986 2058 361222 2294
rect 360986 -582 361222 -346
rect 360986 -902 361222 -666
rect 364686 329758 364922 329994
rect 364686 293758 364922 293994
rect 364686 257758 364922 257994
rect 364686 221758 364922 221994
rect 364686 185758 364922 185994
rect 364686 149758 364922 149994
rect 364686 113758 364922 113994
rect 364686 77758 364922 77994
rect 364686 41758 364922 41994
rect 364686 5758 364922 5994
rect 364686 -2502 364922 -2266
rect 364686 -2822 364922 -2586
rect 372086 337158 372322 337394
rect 368386 333458 368622 333694
rect 368386 297458 368622 297694
rect 368386 261458 368622 261694
rect 368386 225458 368622 225694
rect 368386 189458 368622 189694
rect 368386 153458 368622 153694
rect 368386 117458 368622 117694
rect 368386 81458 368622 81694
rect 368386 45458 368622 45694
rect 368386 9458 368622 9694
rect 368386 -4422 368622 -4186
rect 368386 -4742 368622 -4506
rect 372086 301158 372322 301394
rect 372086 265158 372322 265394
rect 372086 229158 372322 229394
rect 372086 193158 372322 193394
rect 372086 157158 372322 157394
rect 372086 121158 372322 121394
rect 372086 85158 372322 85394
rect 372086 49158 372322 49394
rect 372086 13158 372322 13394
rect 354086 -7302 354322 -7066
rect 354086 -7622 354322 -7386
rect 378986 308058 379222 308294
rect 378986 272058 379222 272294
rect 378986 236058 379222 236294
rect 378986 200058 379222 200294
rect 378986 164058 379222 164294
rect 378986 128058 379222 128294
rect 378986 92058 379222 92294
rect 378986 56058 379222 56294
rect 378986 20058 379222 20294
rect 378986 -1542 379222 -1306
rect 378986 -1862 379222 -1626
rect 382686 311758 382922 311994
rect 382686 275758 382922 275994
rect 382686 239758 382922 239994
rect 382686 203758 382922 203994
rect 382686 167758 382922 167994
rect 382686 131758 382922 131994
rect 382686 95758 382922 95994
rect 382686 59758 382922 59994
rect 382686 23758 382922 23994
rect 382686 -3462 382922 -3226
rect 382686 -3782 382922 -3546
rect 386386 315458 386622 315694
rect 386386 279458 386622 279694
rect 386386 243458 386622 243694
rect 386386 207458 386622 207694
rect 386386 171458 386622 171694
rect 386386 135458 386622 135694
rect 386386 99458 386622 99694
rect 386386 63458 386622 63694
rect 386386 27458 386622 27694
rect 386386 -5382 386622 -5146
rect 386386 -5702 386622 -5466
rect 390086 319158 390322 319394
rect 390086 283158 390322 283394
rect 390086 247158 390322 247394
rect 390086 211158 390322 211394
rect 390086 175158 390322 175394
rect 390086 139158 390322 139394
rect 390086 103158 390322 103394
rect 390086 67158 390322 67394
rect 390086 31158 390322 31394
rect 372086 -6342 372322 -6106
rect 372086 -6662 372322 -6426
rect 396986 326058 397222 326294
rect 396986 290058 397222 290294
rect 396986 254058 397222 254294
rect 396986 218058 397222 218294
rect 396986 182058 397222 182294
rect 396986 146058 397222 146294
rect 396986 110058 397222 110294
rect 396986 74058 397222 74294
rect 396986 38058 397222 38294
rect 396986 2058 397222 2294
rect 396986 -582 397222 -346
rect 396986 -902 397222 -666
rect 400686 329758 400922 329994
rect 400686 293758 400922 293994
rect 400686 257758 400922 257994
rect 400686 221758 400922 221994
rect 400686 185758 400922 185994
rect 400686 149758 400922 149994
rect 400686 113758 400922 113994
rect 400686 77758 400922 77994
rect 400686 41758 400922 41994
rect 400686 5758 400922 5994
rect 400686 -2502 400922 -2266
rect 400686 -2822 400922 -2586
rect 404386 333458 404622 333694
rect 404386 297458 404622 297694
rect 404386 261458 404622 261694
rect 404386 225458 404622 225694
rect 404386 189458 404622 189694
rect 404386 153458 404622 153694
rect 404386 117458 404622 117694
rect 404386 81458 404622 81694
rect 404386 45458 404622 45694
rect 404386 9458 404622 9694
rect 404386 -4422 404622 -4186
rect 404386 -4742 404622 -4506
rect 408086 337158 408322 337394
rect 408086 301158 408322 301394
rect 408086 265158 408322 265394
rect 408086 229158 408322 229394
rect 408086 193158 408322 193394
rect 408086 157158 408322 157394
rect 408086 121158 408322 121394
rect 408086 85158 408322 85394
rect 408086 49158 408322 49394
rect 408086 13158 408322 13394
rect 390086 -7302 390322 -7066
rect 390086 -7622 390322 -7386
rect 414986 308058 415222 308294
rect 414986 272058 415222 272294
rect 414986 236058 415222 236294
rect 414986 200058 415222 200294
rect 414986 164058 415222 164294
rect 414986 128058 415222 128294
rect 414986 92058 415222 92294
rect 414986 56058 415222 56294
rect 414986 20058 415222 20294
rect 414986 -1542 415222 -1306
rect 414986 -1862 415222 -1626
rect 418686 311758 418922 311994
rect 418686 275758 418922 275994
rect 418686 239758 418922 239994
rect 418686 203758 418922 203994
rect 418686 167758 418922 167994
rect 418686 131758 418922 131994
rect 418686 95758 418922 95994
rect 418686 59758 418922 59994
rect 418686 23758 418922 23994
rect 418686 -3462 418922 -3226
rect 418686 -3782 418922 -3546
rect 422386 315458 422622 315694
rect 422386 279458 422622 279694
rect 422386 243458 422622 243694
rect 422386 207458 422622 207694
rect 422386 171458 422622 171694
rect 422386 135458 422622 135694
rect 422386 99458 422622 99694
rect 422386 63458 422622 63694
rect 422386 27458 422622 27694
rect 422386 -5382 422622 -5146
rect 422386 -5702 422622 -5466
rect 426086 319158 426322 319394
rect 426086 283158 426322 283394
rect 426086 247158 426322 247394
rect 426086 211158 426322 211394
rect 426086 175158 426322 175394
rect 426086 139158 426322 139394
rect 426086 103158 426322 103394
rect 426086 67158 426322 67394
rect 426086 31158 426322 31394
rect 408086 -6342 408322 -6106
rect 408086 -6662 408322 -6426
rect 432986 326058 433222 326294
rect 432986 290058 433222 290294
rect 432986 254058 433222 254294
rect 432986 218058 433222 218294
rect 432986 182058 433222 182294
rect 432986 146058 433222 146294
rect 432986 110058 433222 110294
rect 432986 74058 433222 74294
rect 432986 38058 433222 38294
rect 432986 2058 433222 2294
rect 432986 -582 433222 -346
rect 432986 -902 433222 -666
rect 436686 329758 436922 329994
rect 436686 293758 436922 293994
rect 436686 257758 436922 257994
rect 436686 221758 436922 221994
rect 436686 185758 436922 185994
rect 436686 149758 436922 149994
rect 436686 113758 436922 113994
rect 436686 77758 436922 77994
rect 436686 41758 436922 41994
rect 436686 5758 436922 5994
rect 436686 -2502 436922 -2266
rect 436686 -2822 436922 -2586
rect 440386 333458 440622 333694
rect 440386 297458 440622 297694
rect 440386 261458 440622 261694
rect 440386 225458 440622 225694
rect 440386 189458 440622 189694
rect 440386 153458 440622 153694
rect 440386 117458 440622 117694
rect 440386 81458 440622 81694
rect 440386 45458 440622 45694
rect 440386 9458 440622 9694
rect 440386 -4422 440622 -4186
rect 440386 -4742 440622 -4506
rect 444086 337158 444322 337394
rect 444086 301158 444322 301394
rect 444086 265158 444322 265394
rect 444086 229158 444322 229394
rect 444086 193158 444322 193394
rect 444086 157158 444322 157394
rect 444086 121158 444322 121394
rect 444086 85158 444322 85394
rect 444086 49158 444322 49394
rect 444086 13158 444322 13394
rect 426086 -7302 426322 -7066
rect 426086 -7622 426322 -7386
rect 450986 308058 451222 308294
rect 450986 272058 451222 272294
rect 450986 236058 451222 236294
rect 450986 200058 451222 200294
rect 450986 164058 451222 164294
rect 450986 128058 451222 128294
rect 450986 92058 451222 92294
rect 450986 56058 451222 56294
rect 450986 20058 451222 20294
rect 450986 -1542 451222 -1306
rect 450986 -1862 451222 -1626
rect 454686 311758 454922 311994
rect 454686 275758 454922 275994
rect 454686 239758 454922 239994
rect 454686 203758 454922 203994
rect 454686 167758 454922 167994
rect 454686 131758 454922 131994
rect 454686 95758 454922 95994
rect 454686 59758 454922 59994
rect 454686 23758 454922 23994
rect 454686 -3462 454922 -3226
rect 454686 -3782 454922 -3546
rect 458386 315458 458622 315694
rect 458386 279458 458622 279694
rect 458386 243458 458622 243694
rect 458386 207458 458622 207694
rect 458386 171458 458622 171694
rect 458386 135458 458622 135694
rect 458386 99458 458622 99694
rect 458386 63458 458622 63694
rect 458386 27458 458622 27694
rect 458386 -5382 458622 -5146
rect 458386 -5702 458622 -5466
rect 462086 319158 462322 319394
rect 462086 283158 462322 283394
rect 462086 247158 462322 247394
rect 462086 211158 462322 211394
rect 462086 175158 462322 175394
rect 462086 139158 462322 139394
rect 462086 103158 462322 103394
rect 462086 67158 462322 67394
rect 462086 31158 462322 31394
rect 444086 -6342 444322 -6106
rect 444086 -6662 444322 -6426
rect 468986 326058 469222 326294
rect 468986 290058 469222 290294
rect 468986 254058 469222 254294
rect 468986 218058 469222 218294
rect 468986 182058 469222 182294
rect 468986 146058 469222 146294
rect 468986 110058 469222 110294
rect 468986 74058 469222 74294
rect 468986 38058 469222 38294
rect 468986 2058 469222 2294
rect 468986 -582 469222 -346
rect 468986 -902 469222 -666
rect 472686 329758 472922 329994
rect 472686 293758 472922 293994
rect 472686 257758 472922 257994
rect 472686 221758 472922 221994
rect 472686 185758 472922 185994
rect 472686 149758 472922 149994
rect 472686 113758 472922 113994
rect 472686 77758 472922 77994
rect 472686 41758 472922 41994
rect 472686 5758 472922 5994
rect 472686 -2502 472922 -2266
rect 472686 -2822 472922 -2586
rect 476386 333458 476622 333694
rect 476386 297458 476622 297694
rect 476386 261458 476622 261694
rect 476386 225458 476622 225694
rect 476386 189458 476622 189694
rect 476386 153458 476622 153694
rect 476386 117458 476622 117694
rect 476386 81458 476622 81694
rect 476386 45458 476622 45694
rect 476386 9458 476622 9694
rect 476386 -4422 476622 -4186
rect 476386 -4742 476622 -4506
rect 480086 337158 480322 337394
rect 480086 301158 480322 301394
rect 480086 265158 480322 265394
rect 480086 229158 480322 229394
rect 480086 193158 480322 193394
rect 480086 157158 480322 157394
rect 480086 121158 480322 121394
rect 480086 85158 480322 85394
rect 480086 49158 480322 49394
rect 480086 13158 480322 13394
rect 462086 -7302 462322 -7066
rect 462086 -7622 462322 -7386
rect 486986 705562 487222 705798
rect 486986 705242 487222 705478
rect 486986 668058 487222 668294
rect 486986 632058 487222 632294
rect 486986 596058 487222 596294
rect 486986 560058 487222 560294
rect 486986 524058 487222 524294
rect 486986 488058 487222 488294
rect 486986 452058 487222 452294
rect 486986 416058 487222 416294
rect 486986 380058 487222 380294
rect 486986 344058 487222 344294
rect 486986 308058 487222 308294
rect 486986 272058 487222 272294
rect 486986 236058 487222 236294
rect 486986 200058 487222 200294
rect 486986 164058 487222 164294
rect 486986 128058 487222 128294
rect 486986 92058 487222 92294
rect 486986 56058 487222 56294
rect 486986 20058 487222 20294
rect 486986 -1542 487222 -1306
rect 486986 -1862 487222 -1626
rect 490686 671758 490922 671994
rect 490686 635758 490922 635994
rect 490686 599758 490922 599994
rect 490686 563758 490922 563994
rect 490686 527758 490922 527994
rect 490686 491758 490922 491994
rect 490686 455758 490922 455994
rect 490686 419758 490922 419994
rect 490686 383758 490922 383994
rect 490686 347758 490922 347994
rect 490686 311758 490922 311994
rect 490686 275758 490922 275994
rect 490686 239758 490922 239994
rect 490686 203758 490922 203994
rect 490686 167758 490922 167994
rect 490686 131758 490922 131994
rect 490686 95758 490922 95994
rect 490686 59758 490922 59994
rect 490686 23758 490922 23994
rect 490686 -3462 490922 -3226
rect 490686 -3782 490922 -3546
rect 494386 675458 494622 675694
rect 494386 639458 494622 639694
rect 494386 603458 494622 603694
rect 494386 567458 494622 567694
rect 494386 531458 494622 531694
rect 494386 495458 494622 495694
rect 494386 459458 494622 459694
rect 494386 423458 494622 423694
rect 494386 387458 494622 387694
rect 494386 351458 494622 351694
rect 494386 315458 494622 315694
rect 494386 279458 494622 279694
rect 494386 243458 494622 243694
rect 494386 207458 494622 207694
rect 494386 171458 494622 171694
rect 494386 135458 494622 135694
rect 494386 99458 494622 99694
rect 494386 63458 494622 63694
rect 494386 27458 494622 27694
rect 494386 -5382 494622 -5146
rect 494386 -5702 494622 -5466
rect 516086 710362 516322 710598
rect 516086 710042 516322 710278
rect 512386 708442 512622 708678
rect 512386 708122 512622 708358
rect 508686 706522 508922 706758
rect 508686 706202 508922 706438
rect 498086 679158 498322 679394
rect 498086 643158 498322 643394
rect 498086 607158 498322 607394
rect 498086 571158 498322 571394
rect 498086 535158 498322 535394
rect 498086 499158 498322 499394
rect 498086 463158 498322 463394
rect 498086 427158 498322 427394
rect 498086 391158 498322 391394
rect 498086 355158 498322 355394
rect 498086 319158 498322 319394
rect 498086 283158 498322 283394
rect 498086 247158 498322 247394
rect 498086 211158 498322 211394
rect 498086 175158 498322 175394
rect 498086 139158 498322 139394
rect 498086 103158 498322 103394
rect 498086 67158 498322 67394
rect 498086 31158 498322 31394
rect 480086 -6342 480322 -6106
rect 480086 -6662 480322 -6426
rect 504986 704602 505222 704838
rect 504986 704282 505222 704518
rect 504986 686058 505222 686294
rect 504986 650058 505222 650294
rect 504986 614058 505222 614294
rect 504986 578058 505222 578294
rect 504986 542058 505222 542294
rect 504986 506058 505222 506294
rect 504986 470058 505222 470294
rect 504986 434058 505222 434294
rect 504986 398058 505222 398294
rect 504986 362058 505222 362294
rect 504986 326058 505222 326294
rect 504986 290058 505222 290294
rect 504986 254058 505222 254294
rect 504986 218058 505222 218294
rect 504986 182058 505222 182294
rect 504986 146058 505222 146294
rect 504986 110058 505222 110294
rect 504986 74058 505222 74294
rect 504986 38058 505222 38294
rect 504986 2058 505222 2294
rect 504986 -582 505222 -346
rect 504986 -902 505222 -666
rect 508686 689758 508922 689994
rect 508686 653758 508922 653994
rect 508686 617758 508922 617994
rect 508686 581758 508922 581994
rect 508686 545758 508922 545994
rect 508686 509758 508922 509994
rect 508686 473758 508922 473994
rect 508686 437758 508922 437994
rect 508686 401758 508922 401994
rect 508686 365758 508922 365994
rect 508686 329758 508922 329994
rect 508686 293758 508922 293994
rect 508686 257758 508922 257994
rect 508686 221758 508922 221994
rect 508686 185758 508922 185994
rect 508686 149758 508922 149994
rect 508686 113758 508922 113994
rect 508686 77758 508922 77994
rect 508686 41758 508922 41994
rect 508686 5758 508922 5994
rect 508686 -2502 508922 -2266
rect 508686 -2822 508922 -2586
rect 512386 693458 512622 693694
rect 512386 657458 512622 657694
rect 512386 621458 512622 621694
rect 512386 585458 512622 585694
rect 512386 549458 512622 549694
rect 512386 513458 512622 513694
rect 512386 477458 512622 477694
rect 512386 441458 512622 441694
rect 512386 405458 512622 405694
rect 512386 369458 512622 369694
rect 512386 333458 512622 333694
rect 512386 297458 512622 297694
rect 512386 261458 512622 261694
rect 512386 225458 512622 225694
rect 512386 189458 512622 189694
rect 512386 153458 512622 153694
rect 512386 117458 512622 117694
rect 512386 81458 512622 81694
rect 512386 45458 512622 45694
rect 512386 9458 512622 9694
rect 512386 -4422 512622 -4186
rect 512386 -4742 512622 -4506
rect 534086 711322 534322 711558
rect 534086 711002 534322 711238
rect 530386 709402 530622 709638
rect 530386 709082 530622 709318
rect 526686 707482 526922 707718
rect 526686 707162 526922 707398
rect 516086 697158 516322 697394
rect 516086 661158 516322 661394
rect 516086 625158 516322 625394
rect 516086 589158 516322 589394
rect 516086 553158 516322 553394
rect 516086 517158 516322 517394
rect 516086 481158 516322 481394
rect 516086 445158 516322 445394
rect 516086 409158 516322 409394
rect 516086 373158 516322 373394
rect 516086 337158 516322 337394
rect 516086 301158 516322 301394
rect 516086 265158 516322 265394
rect 516086 229158 516322 229394
rect 516086 193158 516322 193394
rect 516086 157158 516322 157394
rect 516086 121158 516322 121394
rect 516086 85158 516322 85394
rect 516086 49158 516322 49394
rect 516086 13158 516322 13394
rect 498086 -7302 498322 -7066
rect 498086 -7622 498322 -7386
rect 522986 705562 523222 705798
rect 522986 705242 523222 705478
rect 522986 668058 523222 668294
rect 522986 632058 523222 632294
rect 522986 596058 523222 596294
rect 522986 560058 523222 560294
rect 522986 524058 523222 524294
rect 522986 488058 523222 488294
rect 522986 452058 523222 452294
rect 522986 416058 523222 416294
rect 522986 380058 523222 380294
rect 522986 344058 523222 344294
rect 522986 308058 523222 308294
rect 522986 272058 523222 272294
rect 522986 236058 523222 236294
rect 522986 200058 523222 200294
rect 522986 164058 523222 164294
rect 522986 128058 523222 128294
rect 522986 92058 523222 92294
rect 522986 56058 523222 56294
rect 522986 20058 523222 20294
rect 522986 -1542 523222 -1306
rect 522986 -1862 523222 -1626
rect 526686 671758 526922 671994
rect 526686 635758 526922 635994
rect 526686 599758 526922 599994
rect 526686 563758 526922 563994
rect 526686 527758 526922 527994
rect 526686 491758 526922 491994
rect 526686 455758 526922 455994
rect 526686 419758 526922 419994
rect 526686 383758 526922 383994
rect 526686 347758 526922 347994
rect 526686 311758 526922 311994
rect 526686 275758 526922 275994
rect 526686 239758 526922 239994
rect 526686 203758 526922 203994
rect 526686 167758 526922 167994
rect 526686 131758 526922 131994
rect 526686 95758 526922 95994
rect 526686 59758 526922 59994
rect 526686 23758 526922 23994
rect 526686 -3462 526922 -3226
rect 526686 -3782 526922 -3546
rect 530386 675458 530622 675694
rect 530386 639458 530622 639694
rect 530386 603458 530622 603694
rect 530386 567458 530622 567694
rect 530386 531458 530622 531694
rect 530386 495458 530622 495694
rect 530386 459458 530622 459694
rect 530386 423458 530622 423694
rect 530386 387458 530622 387694
rect 530386 351458 530622 351694
rect 530386 315458 530622 315694
rect 530386 279458 530622 279694
rect 530386 243458 530622 243694
rect 530386 207458 530622 207694
rect 530386 171458 530622 171694
rect 530386 135458 530622 135694
rect 530386 99458 530622 99694
rect 530386 63458 530622 63694
rect 530386 27458 530622 27694
rect 530386 -5382 530622 -5146
rect 530386 -5702 530622 -5466
rect 552086 710362 552322 710598
rect 552086 710042 552322 710278
rect 548386 708442 548622 708678
rect 548386 708122 548622 708358
rect 544686 706522 544922 706758
rect 544686 706202 544922 706438
rect 534086 679158 534322 679394
rect 534086 643158 534322 643394
rect 534086 607158 534322 607394
rect 534086 571158 534322 571394
rect 534086 535158 534322 535394
rect 534086 499158 534322 499394
rect 534086 463158 534322 463394
rect 534086 427158 534322 427394
rect 534086 391158 534322 391394
rect 534086 355158 534322 355394
rect 534086 319158 534322 319394
rect 534086 283158 534322 283394
rect 534086 247158 534322 247394
rect 534086 211158 534322 211394
rect 534086 175158 534322 175394
rect 534086 139158 534322 139394
rect 534086 103158 534322 103394
rect 534086 67158 534322 67394
rect 534086 31158 534322 31394
rect 516086 -6342 516322 -6106
rect 516086 -6662 516322 -6426
rect 540986 704602 541222 704838
rect 540986 704282 541222 704518
rect 540986 686058 541222 686294
rect 540986 650058 541222 650294
rect 540986 614058 541222 614294
rect 540986 578058 541222 578294
rect 540986 542058 541222 542294
rect 540986 506058 541222 506294
rect 540986 470058 541222 470294
rect 540986 434058 541222 434294
rect 540986 398058 541222 398294
rect 540986 362058 541222 362294
rect 540986 326058 541222 326294
rect 540986 290058 541222 290294
rect 540986 254058 541222 254294
rect 540986 218058 541222 218294
rect 540986 182058 541222 182294
rect 540986 146058 541222 146294
rect 540986 110058 541222 110294
rect 540986 74058 541222 74294
rect 540986 38058 541222 38294
rect 540986 2058 541222 2294
rect 540986 -582 541222 -346
rect 540986 -902 541222 -666
rect 544686 689758 544922 689994
rect 544686 653758 544922 653994
rect 544686 617758 544922 617994
rect 544686 581758 544922 581994
rect 544686 545758 544922 545994
rect 544686 509758 544922 509994
rect 544686 473758 544922 473994
rect 544686 437758 544922 437994
rect 544686 401758 544922 401994
rect 544686 365758 544922 365994
rect 544686 329758 544922 329994
rect 544686 293758 544922 293994
rect 544686 257758 544922 257994
rect 544686 221758 544922 221994
rect 544686 185758 544922 185994
rect 544686 149758 544922 149994
rect 544686 113758 544922 113994
rect 544686 77758 544922 77994
rect 544686 41758 544922 41994
rect 544686 5758 544922 5994
rect 544686 -2502 544922 -2266
rect 544686 -2822 544922 -2586
rect 548386 693458 548622 693694
rect 548386 657458 548622 657694
rect 548386 621458 548622 621694
rect 548386 585458 548622 585694
rect 548386 549458 548622 549694
rect 548386 513458 548622 513694
rect 548386 477458 548622 477694
rect 548386 441458 548622 441694
rect 548386 405458 548622 405694
rect 548386 369458 548622 369694
rect 548386 333458 548622 333694
rect 548386 297458 548622 297694
rect 548386 261458 548622 261694
rect 548386 225458 548622 225694
rect 548386 189458 548622 189694
rect 548386 153458 548622 153694
rect 548386 117458 548622 117694
rect 548386 81458 548622 81694
rect 548386 45458 548622 45694
rect 548386 9458 548622 9694
rect 548386 -4422 548622 -4186
rect 548386 -4742 548622 -4506
rect 570086 711322 570322 711558
rect 570086 711002 570322 711238
rect 566386 709402 566622 709638
rect 566386 709082 566622 709318
rect 562686 707482 562922 707718
rect 562686 707162 562922 707398
rect 552086 697158 552322 697394
rect 552086 661158 552322 661394
rect 552086 625158 552322 625394
rect 552086 589158 552322 589394
rect 552086 553158 552322 553394
rect 552086 517158 552322 517394
rect 552086 481158 552322 481394
rect 552086 445158 552322 445394
rect 552086 409158 552322 409394
rect 552086 373158 552322 373394
rect 552086 337158 552322 337394
rect 552086 301158 552322 301394
rect 552086 265158 552322 265394
rect 552086 229158 552322 229394
rect 552086 193158 552322 193394
rect 552086 157158 552322 157394
rect 552086 121158 552322 121394
rect 552086 85158 552322 85394
rect 552086 49158 552322 49394
rect 552086 13158 552322 13394
rect 534086 -7302 534322 -7066
rect 534086 -7622 534322 -7386
rect 558986 705562 559222 705798
rect 558986 705242 559222 705478
rect 558986 668058 559222 668294
rect 558986 632058 559222 632294
rect 558986 596058 559222 596294
rect 558986 560058 559222 560294
rect 558986 524058 559222 524294
rect 558986 488058 559222 488294
rect 558986 452058 559222 452294
rect 558986 416058 559222 416294
rect 558986 380058 559222 380294
rect 558986 344058 559222 344294
rect 558986 308058 559222 308294
rect 558986 272058 559222 272294
rect 558986 236058 559222 236294
rect 558986 200058 559222 200294
rect 558986 164058 559222 164294
rect 558986 128058 559222 128294
rect 558986 92058 559222 92294
rect 558986 56058 559222 56294
rect 558986 20058 559222 20294
rect 558986 -1542 559222 -1306
rect 558986 -1862 559222 -1626
rect 562686 671758 562922 671994
rect 562686 635758 562922 635994
rect 562686 599758 562922 599994
rect 562686 563758 562922 563994
rect 562686 527758 562922 527994
rect 562686 491758 562922 491994
rect 562686 455758 562922 455994
rect 562686 419758 562922 419994
rect 562686 383758 562922 383994
rect 562686 347758 562922 347994
rect 562686 311758 562922 311994
rect 562686 275758 562922 275994
rect 562686 239758 562922 239994
rect 562686 203758 562922 203994
rect 562686 167758 562922 167994
rect 562686 131758 562922 131994
rect 562686 95758 562922 95994
rect 562686 59758 562922 59994
rect 562686 23758 562922 23994
rect 562686 -3462 562922 -3226
rect 562686 -3782 562922 -3546
rect 566386 675458 566622 675694
rect 566386 639458 566622 639694
rect 566386 603458 566622 603694
rect 566386 567458 566622 567694
rect 566386 531458 566622 531694
rect 566386 495458 566622 495694
rect 566386 459458 566622 459694
rect 566386 423458 566622 423694
rect 566386 387458 566622 387694
rect 566386 351458 566622 351694
rect 566386 315458 566622 315694
rect 566386 279458 566622 279694
rect 566386 243458 566622 243694
rect 566386 207458 566622 207694
rect 566386 171458 566622 171694
rect 566386 135458 566622 135694
rect 566386 99458 566622 99694
rect 566386 63458 566622 63694
rect 566386 27458 566622 27694
rect 566386 -5382 566622 -5146
rect 566386 -5702 566622 -5466
rect 592062 711322 592298 711558
rect 592382 711322 592618 711558
rect 592062 711002 592298 711238
rect 592382 711002 592618 711238
rect 591102 710362 591338 710598
rect 591422 710362 591658 710598
rect 591102 710042 591338 710278
rect 591422 710042 591658 710278
rect 590142 709402 590378 709638
rect 590462 709402 590698 709638
rect 590142 709082 590378 709318
rect 590462 709082 590698 709318
rect 589182 708442 589418 708678
rect 589502 708442 589738 708678
rect 589182 708122 589418 708358
rect 589502 708122 589738 708358
rect 588222 707482 588458 707718
rect 588542 707482 588778 707718
rect 588222 707162 588458 707398
rect 588542 707162 588778 707398
rect 580686 706522 580922 706758
rect 580686 706202 580922 706438
rect 570086 679158 570322 679394
rect 570086 643158 570322 643394
rect 570086 607158 570322 607394
rect 570086 571158 570322 571394
rect 570086 535158 570322 535394
rect 570086 499158 570322 499394
rect 570086 463158 570322 463394
rect 570086 427158 570322 427394
rect 570086 391158 570322 391394
rect 570086 355158 570322 355394
rect 570086 319158 570322 319394
rect 570086 283158 570322 283394
rect 570086 247158 570322 247394
rect 570086 211158 570322 211394
rect 570086 175158 570322 175394
rect 570086 139158 570322 139394
rect 570086 103158 570322 103394
rect 570086 67158 570322 67394
rect 570086 31158 570322 31394
rect 552086 -6342 552322 -6106
rect 552086 -6662 552322 -6426
rect 576986 704602 577222 704838
rect 576986 704282 577222 704518
rect 576986 686058 577222 686294
rect 576986 650058 577222 650294
rect 576986 614058 577222 614294
rect 576986 578058 577222 578294
rect 576986 542058 577222 542294
rect 576986 506058 577222 506294
rect 576986 470058 577222 470294
rect 576986 434058 577222 434294
rect 576986 398058 577222 398294
rect 576986 362058 577222 362294
rect 576986 326058 577222 326294
rect 576986 290058 577222 290294
rect 576986 254058 577222 254294
rect 576986 218058 577222 218294
rect 576986 182058 577222 182294
rect 576986 146058 577222 146294
rect 576986 110058 577222 110294
rect 576986 74058 577222 74294
rect 576986 38058 577222 38294
rect 576986 2058 577222 2294
rect 576986 -582 577222 -346
rect 576986 -902 577222 -666
rect 587262 706522 587498 706758
rect 587582 706522 587818 706758
rect 587262 706202 587498 706438
rect 587582 706202 587818 706438
rect 586302 705562 586538 705798
rect 586622 705562 586858 705798
rect 586302 705242 586538 705478
rect 586622 705242 586858 705478
rect 580686 689758 580922 689994
rect 580686 653758 580922 653994
rect 580686 617758 580922 617994
rect 580686 581758 580922 581994
rect 580686 545758 580922 545994
rect 580686 509758 580922 509994
rect 580686 473758 580922 473994
rect 580686 437758 580922 437994
rect 580686 401758 580922 401994
rect 580686 365758 580922 365994
rect 580686 329758 580922 329994
rect 580686 293758 580922 293994
rect 580686 257758 580922 257994
rect 580686 221758 580922 221994
rect 580686 185758 580922 185994
rect 580686 149758 580922 149994
rect 580686 113758 580922 113994
rect 580686 77758 580922 77994
rect 580686 41758 580922 41994
rect 580686 5758 580922 5994
rect 585342 704602 585578 704838
rect 585662 704602 585898 704838
rect 585342 704282 585578 704518
rect 585662 704282 585898 704518
rect 585342 686058 585578 686294
rect 585662 686058 585898 686294
rect 585342 650058 585578 650294
rect 585662 650058 585898 650294
rect 585342 614058 585578 614294
rect 585662 614058 585898 614294
rect 585342 578058 585578 578294
rect 585662 578058 585898 578294
rect 585342 542058 585578 542294
rect 585662 542058 585898 542294
rect 585342 506058 585578 506294
rect 585662 506058 585898 506294
rect 585342 470058 585578 470294
rect 585662 470058 585898 470294
rect 585342 434058 585578 434294
rect 585662 434058 585898 434294
rect 585342 398058 585578 398294
rect 585662 398058 585898 398294
rect 585342 362058 585578 362294
rect 585662 362058 585898 362294
rect 585342 326058 585578 326294
rect 585662 326058 585898 326294
rect 585342 290058 585578 290294
rect 585662 290058 585898 290294
rect 585342 254058 585578 254294
rect 585662 254058 585898 254294
rect 585342 218058 585578 218294
rect 585662 218058 585898 218294
rect 585342 182058 585578 182294
rect 585662 182058 585898 182294
rect 585342 146058 585578 146294
rect 585662 146058 585898 146294
rect 585342 110058 585578 110294
rect 585662 110058 585898 110294
rect 585342 74058 585578 74294
rect 585662 74058 585898 74294
rect 585342 38058 585578 38294
rect 585662 38058 585898 38294
rect 585342 2058 585578 2294
rect 585662 2058 585898 2294
rect 585342 -582 585578 -346
rect 585662 -582 585898 -346
rect 585342 -902 585578 -666
rect 585662 -902 585898 -666
rect 586302 668058 586538 668294
rect 586622 668058 586858 668294
rect 586302 632058 586538 632294
rect 586622 632058 586858 632294
rect 586302 596058 586538 596294
rect 586622 596058 586858 596294
rect 586302 560058 586538 560294
rect 586622 560058 586858 560294
rect 586302 524058 586538 524294
rect 586622 524058 586858 524294
rect 586302 488058 586538 488294
rect 586622 488058 586858 488294
rect 586302 452058 586538 452294
rect 586622 452058 586858 452294
rect 586302 416058 586538 416294
rect 586622 416058 586858 416294
rect 586302 380058 586538 380294
rect 586622 380058 586858 380294
rect 586302 344058 586538 344294
rect 586622 344058 586858 344294
rect 586302 308058 586538 308294
rect 586622 308058 586858 308294
rect 586302 272058 586538 272294
rect 586622 272058 586858 272294
rect 586302 236058 586538 236294
rect 586622 236058 586858 236294
rect 586302 200058 586538 200294
rect 586622 200058 586858 200294
rect 586302 164058 586538 164294
rect 586622 164058 586858 164294
rect 586302 128058 586538 128294
rect 586622 128058 586858 128294
rect 586302 92058 586538 92294
rect 586622 92058 586858 92294
rect 586302 56058 586538 56294
rect 586622 56058 586858 56294
rect 586302 20058 586538 20294
rect 586622 20058 586858 20294
rect 586302 -1542 586538 -1306
rect 586622 -1542 586858 -1306
rect 586302 -1862 586538 -1626
rect 586622 -1862 586858 -1626
rect 587262 689758 587498 689994
rect 587582 689758 587818 689994
rect 587262 653758 587498 653994
rect 587582 653758 587818 653994
rect 587262 617758 587498 617994
rect 587582 617758 587818 617994
rect 587262 581758 587498 581994
rect 587582 581758 587818 581994
rect 587262 545758 587498 545994
rect 587582 545758 587818 545994
rect 587262 509758 587498 509994
rect 587582 509758 587818 509994
rect 587262 473758 587498 473994
rect 587582 473758 587818 473994
rect 587262 437758 587498 437994
rect 587582 437758 587818 437994
rect 587262 401758 587498 401994
rect 587582 401758 587818 401994
rect 587262 365758 587498 365994
rect 587582 365758 587818 365994
rect 587262 329758 587498 329994
rect 587582 329758 587818 329994
rect 587262 293758 587498 293994
rect 587582 293758 587818 293994
rect 587262 257758 587498 257994
rect 587582 257758 587818 257994
rect 587262 221758 587498 221994
rect 587582 221758 587818 221994
rect 587262 185758 587498 185994
rect 587582 185758 587818 185994
rect 587262 149758 587498 149994
rect 587582 149758 587818 149994
rect 587262 113758 587498 113994
rect 587582 113758 587818 113994
rect 587262 77758 587498 77994
rect 587582 77758 587818 77994
rect 587262 41758 587498 41994
rect 587582 41758 587818 41994
rect 587262 5758 587498 5994
rect 587582 5758 587818 5994
rect 580686 -2502 580922 -2266
rect 580686 -2822 580922 -2586
rect 587262 -2502 587498 -2266
rect 587582 -2502 587818 -2266
rect 587262 -2822 587498 -2586
rect 587582 -2822 587818 -2586
rect 588222 671758 588458 671994
rect 588542 671758 588778 671994
rect 588222 635758 588458 635994
rect 588542 635758 588778 635994
rect 588222 599758 588458 599994
rect 588542 599758 588778 599994
rect 588222 563758 588458 563994
rect 588542 563758 588778 563994
rect 588222 527758 588458 527994
rect 588542 527758 588778 527994
rect 588222 491758 588458 491994
rect 588542 491758 588778 491994
rect 588222 455758 588458 455994
rect 588542 455758 588778 455994
rect 588222 419758 588458 419994
rect 588542 419758 588778 419994
rect 588222 383758 588458 383994
rect 588542 383758 588778 383994
rect 588222 347758 588458 347994
rect 588542 347758 588778 347994
rect 588222 311758 588458 311994
rect 588542 311758 588778 311994
rect 588222 275758 588458 275994
rect 588542 275758 588778 275994
rect 588222 239758 588458 239994
rect 588542 239758 588778 239994
rect 588222 203758 588458 203994
rect 588542 203758 588778 203994
rect 588222 167758 588458 167994
rect 588542 167758 588778 167994
rect 588222 131758 588458 131994
rect 588542 131758 588778 131994
rect 588222 95758 588458 95994
rect 588542 95758 588778 95994
rect 588222 59758 588458 59994
rect 588542 59758 588778 59994
rect 588222 23758 588458 23994
rect 588542 23758 588778 23994
rect 588222 -3462 588458 -3226
rect 588542 -3462 588778 -3226
rect 588222 -3782 588458 -3546
rect 588542 -3782 588778 -3546
rect 589182 693458 589418 693694
rect 589502 693458 589738 693694
rect 589182 657458 589418 657694
rect 589502 657458 589738 657694
rect 589182 621458 589418 621694
rect 589502 621458 589738 621694
rect 589182 585458 589418 585694
rect 589502 585458 589738 585694
rect 589182 549458 589418 549694
rect 589502 549458 589738 549694
rect 589182 513458 589418 513694
rect 589502 513458 589738 513694
rect 589182 477458 589418 477694
rect 589502 477458 589738 477694
rect 589182 441458 589418 441694
rect 589502 441458 589738 441694
rect 589182 405458 589418 405694
rect 589502 405458 589738 405694
rect 589182 369458 589418 369694
rect 589502 369458 589738 369694
rect 589182 333458 589418 333694
rect 589502 333458 589738 333694
rect 589182 297458 589418 297694
rect 589502 297458 589738 297694
rect 589182 261458 589418 261694
rect 589502 261458 589738 261694
rect 589182 225458 589418 225694
rect 589502 225458 589738 225694
rect 589182 189458 589418 189694
rect 589502 189458 589738 189694
rect 589182 153458 589418 153694
rect 589502 153458 589738 153694
rect 589182 117458 589418 117694
rect 589502 117458 589738 117694
rect 589182 81458 589418 81694
rect 589502 81458 589738 81694
rect 589182 45458 589418 45694
rect 589502 45458 589738 45694
rect 589182 9458 589418 9694
rect 589502 9458 589738 9694
rect 589182 -4422 589418 -4186
rect 589502 -4422 589738 -4186
rect 589182 -4742 589418 -4506
rect 589502 -4742 589738 -4506
rect 590142 675458 590378 675694
rect 590462 675458 590698 675694
rect 590142 639458 590378 639694
rect 590462 639458 590698 639694
rect 590142 603458 590378 603694
rect 590462 603458 590698 603694
rect 590142 567458 590378 567694
rect 590462 567458 590698 567694
rect 590142 531458 590378 531694
rect 590462 531458 590698 531694
rect 590142 495458 590378 495694
rect 590462 495458 590698 495694
rect 590142 459458 590378 459694
rect 590462 459458 590698 459694
rect 590142 423458 590378 423694
rect 590462 423458 590698 423694
rect 590142 387458 590378 387694
rect 590462 387458 590698 387694
rect 590142 351458 590378 351694
rect 590462 351458 590698 351694
rect 590142 315458 590378 315694
rect 590462 315458 590698 315694
rect 590142 279458 590378 279694
rect 590462 279458 590698 279694
rect 590142 243458 590378 243694
rect 590462 243458 590698 243694
rect 590142 207458 590378 207694
rect 590462 207458 590698 207694
rect 590142 171458 590378 171694
rect 590462 171458 590698 171694
rect 590142 135458 590378 135694
rect 590462 135458 590698 135694
rect 590142 99458 590378 99694
rect 590462 99458 590698 99694
rect 590142 63458 590378 63694
rect 590462 63458 590698 63694
rect 590142 27458 590378 27694
rect 590462 27458 590698 27694
rect 590142 -5382 590378 -5146
rect 590462 -5382 590698 -5146
rect 590142 -5702 590378 -5466
rect 590462 -5702 590698 -5466
rect 591102 697158 591338 697394
rect 591422 697158 591658 697394
rect 591102 661158 591338 661394
rect 591422 661158 591658 661394
rect 591102 625158 591338 625394
rect 591422 625158 591658 625394
rect 591102 589158 591338 589394
rect 591422 589158 591658 589394
rect 591102 553158 591338 553394
rect 591422 553158 591658 553394
rect 591102 517158 591338 517394
rect 591422 517158 591658 517394
rect 591102 481158 591338 481394
rect 591422 481158 591658 481394
rect 591102 445158 591338 445394
rect 591422 445158 591658 445394
rect 591102 409158 591338 409394
rect 591422 409158 591658 409394
rect 591102 373158 591338 373394
rect 591422 373158 591658 373394
rect 591102 337158 591338 337394
rect 591422 337158 591658 337394
rect 591102 301158 591338 301394
rect 591422 301158 591658 301394
rect 591102 265158 591338 265394
rect 591422 265158 591658 265394
rect 591102 229158 591338 229394
rect 591422 229158 591658 229394
rect 591102 193158 591338 193394
rect 591422 193158 591658 193394
rect 591102 157158 591338 157394
rect 591422 157158 591658 157394
rect 591102 121158 591338 121394
rect 591422 121158 591658 121394
rect 591102 85158 591338 85394
rect 591422 85158 591658 85394
rect 591102 49158 591338 49394
rect 591422 49158 591658 49394
rect 591102 13158 591338 13394
rect 591422 13158 591658 13394
rect 591102 -6342 591338 -6106
rect 591422 -6342 591658 -6106
rect 591102 -6662 591338 -6426
rect 591422 -6662 591658 -6426
rect 592062 679158 592298 679394
rect 592382 679158 592618 679394
rect 592062 643158 592298 643394
rect 592382 643158 592618 643394
rect 592062 607158 592298 607394
rect 592382 607158 592618 607394
rect 592062 571158 592298 571394
rect 592382 571158 592618 571394
rect 592062 535158 592298 535394
rect 592382 535158 592618 535394
rect 592062 499158 592298 499394
rect 592382 499158 592618 499394
rect 592062 463158 592298 463394
rect 592382 463158 592618 463394
rect 592062 427158 592298 427394
rect 592382 427158 592618 427394
rect 592062 391158 592298 391394
rect 592382 391158 592618 391394
rect 592062 355158 592298 355394
rect 592382 355158 592618 355394
rect 592062 319158 592298 319394
rect 592382 319158 592618 319394
rect 592062 283158 592298 283394
rect 592382 283158 592618 283394
rect 592062 247158 592298 247394
rect 592382 247158 592618 247394
rect 592062 211158 592298 211394
rect 592382 211158 592618 211394
rect 592062 175158 592298 175394
rect 592382 175158 592618 175394
rect 592062 139158 592298 139394
rect 592382 139158 592618 139394
rect 592062 103158 592298 103394
rect 592382 103158 592618 103394
rect 592062 67158 592298 67394
rect 592382 67158 592618 67394
rect 592062 31158 592298 31394
rect 592382 31158 592618 31394
rect 570086 -7302 570322 -7066
rect 570086 -7622 570322 -7386
rect 592062 -7302 592298 -7066
rect 592382 -7302 592618 -7066
rect 592062 -7622 592298 -7386
rect 592382 -7622 592618 -7386
<< metal5 >>
rect -8726 711558 592650 711590
rect -8726 711322 -8694 711558
rect -8458 711322 -8374 711558
rect -8138 711322 30086 711558
rect 30322 711322 66086 711558
rect 66322 711322 102086 711558
rect 102322 711322 138086 711558
rect 138322 711322 174086 711558
rect 174322 711322 210086 711558
rect 210322 711322 246086 711558
rect 246322 711322 282086 711558
rect 282322 711322 318086 711558
rect 318322 711322 354086 711558
rect 354322 711322 390086 711558
rect 390322 711322 426086 711558
rect 426322 711322 462086 711558
rect 462322 711322 498086 711558
rect 498322 711322 534086 711558
rect 534322 711322 570086 711558
rect 570322 711322 592062 711558
rect 592298 711322 592382 711558
rect 592618 711322 592650 711558
rect -8726 711238 592650 711322
rect -8726 711002 -8694 711238
rect -8458 711002 -8374 711238
rect -8138 711002 30086 711238
rect 30322 711002 66086 711238
rect 66322 711002 102086 711238
rect 102322 711002 138086 711238
rect 138322 711002 174086 711238
rect 174322 711002 210086 711238
rect 210322 711002 246086 711238
rect 246322 711002 282086 711238
rect 282322 711002 318086 711238
rect 318322 711002 354086 711238
rect 354322 711002 390086 711238
rect 390322 711002 426086 711238
rect 426322 711002 462086 711238
rect 462322 711002 498086 711238
rect 498322 711002 534086 711238
rect 534322 711002 570086 711238
rect 570322 711002 592062 711238
rect 592298 711002 592382 711238
rect 592618 711002 592650 711238
rect -8726 710970 592650 711002
rect -7766 710598 591690 710630
rect -7766 710362 -7734 710598
rect -7498 710362 -7414 710598
rect -7178 710362 12086 710598
rect 12322 710362 48086 710598
rect 48322 710362 84086 710598
rect 84322 710362 120086 710598
rect 120322 710362 156086 710598
rect 156322 710362 192086 710598
rect 192322 710362 228086 710598
rect 228322 710362 264086 710598
rect 264322 710362 300086 710598
rect 300322 710362 336086 710598
rect 336322 710362 372086 710598
rect 372322 710362 408086 710598
rect 408322 710362 444086 710598
rect 444322 710362 480086 710598
rect 480322 710362 516086 710598
rect 516322 710362 552086 710598
rect 552322 710362 591102 710598
rect 591338 710362 591422 710598
rect 591658 710362 591690 710598
rect -7766 710278 591690 710362
rect -7766 710042 -7734 710278
rect -7498 710042 -7414 710278
rect -7178 710042 12086 710278
rect 12322 710042 48086 710278
rect 48322 710042 84086 710278
rect 84322 710042 120086 710278
rect 120322 710042 156086 710278
rect 156322 710042 192086 710278
rect 192322 710042 228086 710278
rect 228322 710042 264086 710278
rect 264322 710042 300086 710278
rect 300322 710042 336086 710278
rect 336322 710042 372086 710278
rect 372322 710042 408086 710278
rect 408322 710042 444086 710278
rect 444322 710042 480086 710278
rect 480322 710042 516086 710278
rect 516322 710042 552086 710278
rect 552322 710042 591102 710278
rect 591338 710042 591422 710278
rect 591658 710042 591690 710278
rect -7766 710010 591690 710042
rect -6806 709638 590730 709670
rect -6806 709402 -6774 709638
rect -6538 709402 -6454 709638
rect -6218 709402 26386 709638
rect 26622 709402 62386 709638
rect 62622 709402 98386 709638
rect 98622 709402 134386 709638
rect 134622 709402 170386 709638
rect 170622 709402 206386 709638
rect 206622 709402 242386 709638
rect 242622 709402 278386 709638
rect 278622 709402 314386 709638
rect 314622 709402 350386 709638
rect 350622 709402 386386 709638
rect 386622 709402 422386 709638
rect 422622 709402 458386 709638
rect 458622 709402 494386 709638
rect 494622 709402 530386 709638
rect 530622 709402 566386 709638
rect 566622 709402 590142 709638
rect 590378 709402 590462 709638
rect 590698 709402 590730 709638
rect -6806 709318 590730 709402
rect -6806 709082 -6774 709318
rect -6538 709082 -6454 709318
rect -6218 709082 26386 709318
rect 26622 709082 62386 709318
rect 62622 709082 98386 709318
rect 98622 709082 134386 709318
rect 134622 709082 170386 709318
rect 170622 709082 206386 709318
rect 206622 709082 242386 709318
rect 242622 709082 278386 709318
rect 278622 709082 314386 709318
rect 314622 709082 350386 709318
rect 350622 709082 386386 709318
rect 386622 709082 422386 709318
rect 422622 709082 458386 709318
rect 458622 709082 494386 709318
rect 494622 709082 530386 709318
rect 530622 709082 566386 709318
rect 566622 709082 590142 709318
rect 590378 709082 590462 709318
rect 590698 709082 590730 709318
rect -6806 709050 590730 709082
rect -5846 708678 589770 708710
rect -5846 708442 -5814 708678
rect -5578 708442 -5494 708678
rect -5258 708442 8386 708678
rect 8622 708442 44386 708678
rect 44622 708442 80386 708678
rect 80622 708442 116386 708678
rect 116622 708442 152386 708678
rect 152622 708442 188386 708678
rect 188622 708442 224386 708678
rect 224622 708442 260386 708678
rect 260622 708442 296386 708678
rect 296622 708442 332386 708678
rect 332622 708442 368386 708678
rect 368622 708442 404386 708678
rect 404622 708442 440386 708678
rect 440622 708442 476386 708678
rect 476622 708442 512386 708678
rect 512622 708442 548386 708678
rect 548622 708442 589182 708678
rect 589418 708442 589502 708678
rect 589738 708442 589770 708678
rect -5846 708358 589770 708442
rect -5846 708122 -5814 708358
rect -5578 708122 -5494 708358
rect -5258 708122 8386 708358
rect 8622 708122 44386 708358
rect 44622 708122 80386 708358
rect 80622 708122 116386 708358
rect 116622 708122 152386 708358
rect 152622 708122 188386 708358
rect 188622 708122 224386 708358
rect 224622 708122 260386 708358
rect 260622 708122 296386 708358
rect 296622 708122 332386 708358
rect 332622 708122 368386 708358
rect 368622 708122 404386 708358
rect 404622 708122 440386 708358
rect 440622 708122 476386 708358
rect 476622 708122 512386 708358
rect 512622 708122 548386 708358
rect 548622 708122 589182 708358
rect 589418 708122 589502 708358
rect 589738 708122 589770 708358
rect -5846 708090 589770 708122
rect -4886 707718 588810 707750
rect -4886 707482 -4854 707718
rect -4618 707482 -4534 707718
rect -4298 707482 22686 707718
rect 22922 707482 58686 707718
rect 58922 707482 94686 707718
rect 94922 707482 130686 707718
rect 130922 707482 166686 707718
rect 166922 707482 202686 707718
rect 202922 707482 238686 707718
rect 238922 707482 274686 707718
rect 274922 707482 310686 707718
rect 310922 707482 346686 707718
rect 346922 707482 382686 707718
rect 382922 707482 418686 707718
rect 418922 707482 454686 707718
rect 454922 707482 490686 707718
rect 490922 707482 526686 707718
rect 526922 707482 562686 707718
rect 562922 707482 588222 707718
rect 588458 707482 588542 707718
rect 588778 707482 588810 707718
rect -4886 707398 588810 707482
rect -4886 707162 -4854 707398
rect -4618 707162 -4534 707398
rect -4298 707162 22686 707398
rect 22922 707162 58686 707398
rect 58922 707162 94686 707398
rect 94922 707162 130686 707398
rect 130922 707162 166686 707398
rect 166922 707162 202686 707398
rect 202922 707162 238686 707398
rect 238922 707162 274686 707398
rect 274922 707162 310686 707398
rect 310922 707162 346686 707398
rect 346922 707162 382686 707398
rect 382922 707162 418686 707398
rect 418922 707162 454686 707398
rect 454922 707162 490686 707398
rect 490922 707162 526686 707398
rect 526922 707162 562686 707398
rect 562922 707162 588222 707398
rect 588458 707162 588542 707398
rect 588778 707162 588810 707398
rect -4886 707130 588810 707162
rect -3926 706758 587850 706790
rect -3926 706522 -3894 706758
rect -3658 706522 -3574 706758
rect -3338 706522 4686 706758
rect 4922 706522 40686 706758
rect 40922 706522 76686 706758
rect 76922 706522 112686 706758
rect 112922 706522 148686 706758
rect 148922 706522 184686 706758
rect 184922 706522 220686 706758
rect 220922 706522 256686 706758
rect 256922 706522 292686 706758
rect 292922 706522 328686 706758
rect 328922 706522 364686 706758
rect 364922 706522 400686 706758
rect 400922 706522 436686 706758
rect 436922 706522 472686 706758
rect 472922 706522 508686 706758
rect 508922 706522 544686 706758
rect 544922 706522 580686 706758
rect 580922 706522 587262 706758
rect 587498 706522 587582 706758
rect 587818 706522 587850 706758
rect -3926 706438 587850 706522
rect -3926 706202 -3894 706438
rect -3658 706202 -3574 706438
rect -3338 706202 4686 706438
rect 4922 706202 40686 706438
rect 40922 706202 76686 706438
rect 76922 706202 112686 706438
rect 112922 706202 148686 706438
rect 148922 706202 184686 706438
rect 184922 706202 220686 706438
rect 220922 706202 256686 706438
rect 256922 706202 292686 706438
rect 292922 706202 328686 706438
rect 328922 706202 364686 706438
rect 364922 706202 400686 706438
rect 400922 706202 436686 706438
rect 436922 706202 472686 706438
rect 472922 706202 508686 706438
rect 508922 706202 544686 706438
rect 544922 706202 580686 706438
rect 580922 706202 587262 706438
rect 587498 706202 587582 706438
rect 587818 706202 587850 706438
rect -3926 706170 587850 706202
rect -2966 705798 586890 705830
rect -2966 705562 -2934 705798
rect -2698 705562 -2614 705798
rect -2378 705562 18986 705798
rect 19222 705562 54986 705798
rect 55222 705562 90986 705798
rect 91222 705562 126986 705798
rect 127222 705562 162986 705798
rect 163222 705562 198986 705798
rect 199222 705562 234986 705798
rect 235222 705562 270986 705798
rect 271222 705562 306986 705798
rect 307222 705562 342986 705798
rect 343222 705562 378986 705798
rect 379222 705562 414986 705798
rect 415222 705562 450986 705798
rect 451222 705562 486986 705798
rect 487222 705562 522986 705798
rect 523222 705562 558986 705798
rect 559222 705562 586302 705798
rect 586538 705562 586622 705798
rect 586858 705562 586890 705798
rect -2966 705478 586890 705562
rect -2966 705242 -2934 705478
rect -2698 705242 -2614 705478
rect -2378 705242 18986 705478
rect 19222 705242 54986 705478
rect 55222 705242 90986 705478
rect 91222 705242 126986 705478
rect 127222 705242 162986 705478
rect 163222 705242 198986 705478
rect 199222 705242 234986 705478
rect 235222 705242 270986 705478
rect 271222 705242 306986 705478
rect 307222 705242 342986 705478
rect 343222 705242 378986 705478
rect 379222 705242 414986 705478
rect 415222 705242 450986 705478
rect 451222 705242 486986 705478
rect 487222 705242 522986 705478
rect 523222 705242 558986 705478
rect 559222 705242 586302 705478
rect 586538 705242 586622 705478
rect 586858 705242 586890 705478
rect -2966 705210 586890 705242
rect -2006 704838 585930 704870
rect -2006 704602 -1974 704838
rect -1738 704602 -1654 704838
rect -1418 704602 986 704838
rect 1222 704602 36986 704838
rect 37222 704602 72986 704838
rect 73222 704602 108986 704838
rect 109222 704602 144986 704838
rect 145222 704602 180986 704838
rect 181222 704602 216986 704838
rect 217222 704602 252986 704838
rect 253222 704602 288986 704838
rect 289222 704602 324986 704838
rect 325222 704602 360986 704838
rect 361222 704602 396986 704838
rect 397222 704602 432986 704838
rect 433222 704602 468986 704838
rect 469222 704602 504986 704838
rect 505222 704602 540986 704838
rect 541222 704602 576986 704838
rect 577222 704602 585342 704838
rect 585578 704602 585662 704838
rect 585898 704602 585930 704838
rect -2006 704518 585930 704602
rect -2006 704282 -1974 704518
rect -1738 704282 -1654 704518
rect -1418 704282 986 704518
rect 1222 704282 36986 704518
rect 37222 704282 72986 704518
rect 73222 704282 108986 704518
rect 109222 704282 144986 704518
rect 145222 704282 180986 704518
rect 181222 704282 216986 704518
rect 217222 704282 252986 704518
rect 253222 704282 288986 704518
rect 289222 704282 324986 704518
rect 325222 704282 360986 704518
rect 361222 704282 396986 704518
rect 397222 704282 432986 704518
rect 433222 704282 468986 704518
rect 469222 704282 504986 704518
rect 505222 704282 540986 704518
rect 541222 704282 576986 704518
rect 577222 704282 585342 704518
rect 585578 704282 585662 704518
rect 585898 704282 585930 704518
rect -2006 704250 585930 704282
rect -8726 697394 592650 697576
rect -8726 697158 -7734 697394
rect -7498 697158 -7414 697394
rect -7178 697158 12086 697394
rect 12322 697158 48086 697394
rect 48322 697158 84086 697394
rect 84322 697158 120086 697394
rect 120322 697158 156086 697394
rect 156322 697158 192086 697394
rect 192322 697158 228086 697394
rect 228322 697158 264086 697394
rect 264322 697158 300086 697394
rect 300322 697158 336086 697394
rect 336322 697158 372086 697394
rect 372322 697158 408086 697394
rect 408322 697158 444086 697394
rect 444322 697158 480086 697394
rect 480322 697158 516086 697394
rect 516322 697158 552086 697394
rect 552322 697158 591102 697394
rect 591338 697158 591422 697394
rect 591658 697158 592650 697394
rect -8726 696976 592650 697158
rect -6806 693694 590730 693876
rect -6806 693458 -5814 693694
rect -5578 693458 -5494 693694
rect -5258 693458 8386 693694
rect 8622 693458 44386 693694
rect 44622 693458 80386 693694
rect 80622 693458 116386 693694
rect 116622 693458 152386 693694
rect 152622 693458 188386 693694
rect 188622 693458 224386 693694
rect 224622 693458 260386 693694
rect 260622 693458 296386 693694
rect 296622 693458 332386 693694
rect 332622 693458 368386 693694
rect 368622 693458 404386 693694
rect 404622 693458 440386 693694
rect 440622 693458 476386 693694
rect 476622 693458 512386 693694
rect 512622 693458 548386 693694
rect 548622 693458 589182 693694
rect 589418 693458 589502 693694
rect 589738 693458 590730 693694
rect -6806 693276 590730 693458
rect -4886 689994 588810 690176
rect -4886 689758 -3894 689994
rect -3658 689758 -3574 689994
rect -3338 689758 4686 689994
rect 4922 689758 40686 689994
rect 40922 689758 76686 689994
rect 76922 689758 112686 689994
rect 112922 689758 148686 689994
rect 148922 689758 184686 689994
rect 184922 689758 220686 689994
rect 220922 689758 256686 689994
rect 256922 689758 292686 689994
rect 292922 689758 328686 689994
rect 328922 689758 364686 689994
rect 364922 689758 400686 689994
rect 400922 689758 436686 689994
rect 436922 689758 472686 689994
rect 472922 689758 508686 689994
rect 508922 689758 544686 689994
rect 544922 689758 580686 689994
rect 580922 689758 587262 689994
rect 587498 689758 587582 689994
rect 587818 689758 588810 689994
rect -4886 689576 588810 689758
rect -2966 686294 586890 686476
rect -2966 686058 -1974 686294
rect -1738 686058 -1654 686294
rect -1418 686058 986 686294
rect 1222 686058 36986 686294
rect 37222 686058 72986 686294
rect 73222 686058 108986 686294
rect 109222 686058 144986 686294
rect 145222 686058 180986 686294
rect 181222 686058 216986 686294
rect 217222 686058 252986 686294
rect 253222 686058 288986 686294
rect 289222 686058 324986 686294
rect 325222 686058 360986 686294
rect 361222 686058 396986 686294
rect 397222 686058 432986 686294
rect 433222 686058 468986 686294
rect 469222 686058 504986 686294
rect 505222 686058 540986 686294
rect 541222 686058 576986 686294
rect 577222 686058 585342 686294
rect 585578 686058 585662 686294
rect 585898 686058 586890 686294
rect -2966 685876 586890 686058
rect -8726 679394 592650 679576
rect -8726 679158 -8694 679394
rect -8458 679158 -8374 679394
rect -8138 679158 30086 679394
rect 30322 679158 66086 679394
rect 66322 679158 102086 679394
rect 102322 679158 138086 679394
rect 138322 679158 174086 679394
rect 174322 679158 210086 679394
rect 210322 679158 246086 679394
rect 246322 679158 282086 679394
rect 282322 679158 318086 679394
rect 318322 679158 354086 679394
rect 354322 679158 390086 679394
rect 390322 679158 426086 679394
rect 426322 679158 462086 679394
rect 462322 679158 498086 679394
rect 498322 679158 534086 679394
rect 534322 679158 570086 679394
rect 570322 679158 592062 679394
rect 592298 679158 592382 679394
rect 592618 679158 592650 679394
rect -8726 678976 592650 679158
rect -6806 675694 590730 675876
rect -6806 675458 -6774 675694
rect -6538 675458 -6454 675694
rect -6218 675458 26386 675694
rect 26622 675458 62386 675694
rect 62622 675458 98386 675694
rect 98622 675458 134386 675694
rect 134622 675458 170386 675694
rect 170622 675458 206386 675694
rect 206622 675458 242386 675694
rect 242622 675458 278386 675694
rect 278622 675458 314386 675694
rect 314622 675458 350386 675694
rect 350622 675458 386386 675694
rect 386622 675458 422386 675694
rect 422622 675458 458386 675694
rect 458622 675458 494386 675694
rect 494622 675458 530386 675694
rect 530622 675458 566386 675694
rect 566622 675458 590142 675694
rect 590378 675458 590462 675694
rect 590698 675458 590730 675694
rect -6806 675276 590730 675458
rect -4886 671994 588810 672176
rect -4886 671758 -4854 671994
rect -4618 671758 -4534 671994
rect -4298 671758 22686 671994
rect 22922 671758 58686 671994
rect 58922 671758 94686 671994
rect 94922 671758 130686 671994
rect 130922 671758 166686 671994
rect 166922 671758 202686 671994
rect 202922 671758 238686 671994
rect 238922 671758 274686 671994
rect 274922 671758 310686 671994
rect 310922 671758 346686 671994
rect 346922 671758 382686 671994
rect 382922 671758 418686 671994
rect 418922 671758 454686 671994
rect 454922 671758 490686 671994
rect 490922 671758 526686 671994
rect 526922 671758 562686 671994
rect 562922 671758 588222 671994
rect 588458 671758 588542 671994
rect 588778 671758 588810 671994
rect -4886 671576 588810 671758
rect -2966 668294 586890 668476
rect -2966 668058 -2934 668294
rect -2698 668058 -2614 668294
rect -2378 668058 18986 668294
rect 19222 668058 54986 668294
rect 55222 668058 90986 668294
rect 91222 668058 126986 668294
rect 127222 668058 162986 668294
rect 163222 668058 198986 668294
rect 199222 668058 234986 668294
rect 235222 668058 270986 668294
rect 271222 668058 306986 668294
rect 307222 668058 342986 668294
rect 343222 668058 378986 668294
rect 379222 668058 414986 668294
rect 415222 668058 450986 668294
rect 451222 668058 486986 668294
rect 487222 668058 522986 668294
rect 523222 668058 558986 668294
rect 559222 668058 586302 668294
rect 586538 668058 586622 668294
rect 586858 668058 586890 668294
rect -2966 667876 586890 668058
rect -8726 661394 592650 661576
rect -8726 661158 -7734 661394
rect -7498 661158 -7414 661394
rect -7178 661158 12086 661394
rect 12322 661158 48086 661394
rect 48322 661158 84086 661394
rect 84322 661158 120086 661394
rect 120322 661158 156086 661394
rect 156322 661158 192086 661394
rect 192322 661158 228086 661394
rect 228322 661158 264086 661394
rect 264322 661158 300086 661394
rect 300322 661158 336086 661394
rect 336322 661158 372086 661394
rect 372322 661158 408086 661394
rect 408322 661158 444086 661394
rect 444322 661158 480086 661394
rect 480322 661158 516086 661394
rect 516322 661158 552086 661394
rect 552322 661158 591102 661394
rect 591338 661158 591422 661394
rect 591658 661158 592650 661394
rect -8726 660976 592650 661158
rect -6806 657694 590730 657876
rect -6806 657458 -5814 657694
rect -5578 657458 -5494 657694
rect -5258 657458 8386 657694
rect 8622 657458 44386 657694
rect 44622 657458 80386 657694
rect 80622 657458 116386 657694
rect 116622 657458 152386 657694
rect 152622 657458 188386 657694
rect 188622 657458 224386 657694
rect 224622 657458 260386 657694
rect 260622 657458 296386 657694
rect 296622 657458 332386 657694
rect 332622 657458 368386 657694
rect 368622 657458 404386 657694
rect 404622 657458 440386 657694
rect 440622 657458 476386 657694
rect 476622 657458 512386 657694
rect 512622 657458 548386 657694
rect 548622 657458 589182 657694
rect 589418 657458 589502 657694
rect 589738 657458 590730 657694
rect -6806 657276 590730 657458
rect -4886 653994 588810 654176
rect -4886 653758 -3894 653994
rect -3658 653758 -3574 653994
rect -3338 653758 4686 653994
rect 4922 653758 40686 653994
rect 40922 653758 76686 653994
rect 76922 653758 112686 653994
rect 112922 653758 148686 653994
rect 148922 653758 184686 653994
rect 184922 653758 220686 653994
rect 220922 653758 256686 653994
rect 256922 653758 292686 653994
rect 292922 653758 328686 653994
rect 328922 653758 364686 653994
rect 364922 653758 400686 653994
rect 400922 653758 436686 653994
rect 436922 653758 472686 653994
rect 472922 653758 508686 653994
rect 508922 653758 544686 653994
rect 544922 653758 580686 653994
rect 580922 653758 587262 653994
rect 587498 653758 587582 653994
rect 587818 653758 588810 653994
rect -4886 653576 588810 653758
rect -2966 650294 586890 650476
rect -2966 650058 -1974 650294
rect -1738 650058 -1654 650294
rect -1418 650058 986 650294
rect 1222 650058 36986 650294
rect 37222 650058 72986 650294
rect 73222 650058 108986 650294
rect 109222 650058 144986 650294
rect 145222 650058 180986 650294
rect 181222 650058 216986 650294
rect 217222 650058 252986 650294
rect 253222 650058 288986 650294
rect 289222 650058 324986 650294
rect 325222 650058 360986 650294
rect 361222 650058 396986 650294
rect 397222 650058 432986 650294
rect 433222 650058 468986 650294
rect 469222 650058 504986 650294
rect 505222 650058 540986 650294
rect 541222 650058 576986 650294
rect 577222 650058 585342 650294
rect 585578 650058 585662 650294
rect 585898 650058 586890 650294
rect -2966 649876 586890 650058
rect -8726 643394 592650 643576
rect -8726 643158 -8694 643394
rect -8458 643158 -8374 643394
rect -8138 643158 30086 643394
rect 30322 643158 66086 643394
rect 66322 643158 102086 643394
rect 102322 643158 138086 643394
rect 138322 643158 174086 643394
rect 174322 643158 210086 643394
rect 210322 643158 246086 643394
rect 246322 643158 282086 643394
rect 282322 643158 318086 643394
rect 318322 643158 354086 643394
rect 354322 643158 390086 643394
rect 390322 643158 426086 643394
rect 426322 643158 462086 643394
rect 462322 643158 498086 643394
rect 498322 643158 534086 643394
rect 534322 643158 570086 643394
rect 570322 643158 592062 643394
rect 592298 643158 592382 643394
rect 592618 643158 592650 643394
rect -8726 642976 592650 643158
rect -6806 639694 590730 639876
rect -6806 639458 -6774 639694
rect -6538 639458 -6454 639694
rect -6218 639458 26386 639694
rect 26622 639458 62386 639694
rect 62622 639458 98386 639694
rect 98622 639458 134386 639694
rect 134622 639458 170386 639694
rect 170622 639458 206386 639694
rect 206622 639458 242386 639694
rect 242622 639458 278386 639694
rect 278622 639458 314386 639694
rect 314622 639458 350386 639694
rect 350622 639458 386386 639694
rect 386622 639458 422386 639694
rect 422622 639458 458386 639694
rect 458622 639458 494386 639694
rect 494622 639458 530386 639694
rect 530622 639458 566386 639694
rect 566622 639458 590142 639694
rect 590378 639458 590462 639694
rect 590698 639458 590730 639694
rect -6806 639276 590730 639458
rect -4886 635994 588810 636176
rect -4886 635758 -4854 635994
rect -4618 635758 -4534 635994
rect -4298 635758 22686 635994
rect 22922 635758 58686 635994
rect 58922 635758 94686 635994
rect 94922 635758 130686 635994
rect 130922 635758 166686 635994
rect 166922 635758 202686 635994
rect 202922 635758 238686 635994
rect 238922 635758 274686 635994
rect 274922 635758 310686 635994
rect 310922 635758 346686 635994
rect 346922 635758 382686 635994
rect 382922 635758 418686 635994
rect 418922 635758 454686 635994
rect 454922 635758 490686 635994
rect 490922 635758 526686 635994
rect 526922 635758 562686 635994
rect 562922 635758 588222 635994
rect 588458 635758 588542 635994
rect 588778 635758 588810 635994
rect -4886 635576 588810 635758
rect -2966 632294 586890 632476
rect -2966 632058 -2934 632294
rect -2698 632058 -2614 632294
rect -2378 632058 18986 632294
rect 19222 632058 54986 632294
rect 55222 632058 90986 632294
rect 91222 632058 126986 632294
rect 127222 632058 162986 632294
rect 163222 632058 198986 632294
rect 199222 632058 234986 632294
rect 235222 632058 270986 632294
rect 271222 632058 306986 632294
rect 307222 632058 342986 632294
rect 343222 632058 378986 632294
rect 379222 632058 414986 632294
rect 415222 632058 450986 632294
rect 451222 632058 486986 632294
rect 487222 632058 522986 632294
rect 523222 632058 558986 632294
rect 559222 632058 586302 632294
rect 586538 632058 586622 632294
rect 586858 632058 586890 632294
rect -2966 631876 586890 632058
rect -8726 625394 592650 625576
rect -8726 625158 -7734 625394
rect -7498 625158 -7414 625394
rect -7178 625158 12086 625394
rect 12322 625158 48086 625394
rect 48322 625158 84086 625394
rect 84322 625158 120086 625394
rect 120322 625158 156086 625394
rect 156322 625158 192086 625394
rect 192322 625158 228086 625394
rect 228322 625158 264086 625394
rect 264322 625158 300086 625394
rect 300322 625158 336086 625394
rect 336322 625158 372086 625394
rect 372322 625158 408086 625394
rect 408322 625158 444086 625394
rect 444322 625158 480086 625394
rect 480322 625158 516086 625394
rect 516322 625158 552086 625394
rect 552322 625158 591102 625394
rect 591338 625158 591422 625394
rect 591658 625158 592650 625394
rect -8726 624976 592650 625158
rect -6806 621694 590730 621876
rect -6806 621458 -5814 621694
rect -5578 621458 -5494 621694
rect -5258 621458 8386 621694
rect 8622 621458 44386 621694
rect 44622 621458 80386 621694
rect 80622 621458 116386 621694
rect 116622 621458 152386 621694
rect 152622 621458 188386 621694
rect 188622 621458 224386 621694
rect 224622 621458 260386 621694
rect 260622 621458 296386 621694
rect 296622 621458 332386 621694
rect 332622 621458 368386 621694
rect 368622 621458 404386 621694
rect 404622 621458 440386 621694
rect 440622 621458 476386 621694
rect 476622 621458 512386 621694
rect 512622 621458 548386 621694
rect 548622 621458 589182 621694
rect 589418 621458 589502 621694
rect 589738 621458 590730 621694
rect -6806 621276 590730 621458
rect -4886 617994 588810 618176
rect -4886 617758 -3894 617994
rect -3658 617758 -3574 617994
rect -3338 617758 4686 617994
rect 4922 617758 40686 617994
rect 40922 617758 76686 617994
rect 76922 617758 112686 617994
rect 112922 617758 148686 617994
rect 148922 617758 184686 617994
rect 184922 617758 220686 617994
rect 220922 617758 256686 617994
rect 256922 617758 292686 617994
rect 292922 617758 328686 617994
rect 328922 617758 364686 617994
rect 364922 617758 400686 617994
rect 400922 617758 436686 617994
rect 436922 617758 472686 617994
rect 472922 617758 508686 617994
rect 508922 617758 544686 617994
rect 544922 617758 580686 617994
rect 580922 617758 587262 617994
rect 587498 617758 587582 617994
rect 587818 617758 588810 617994
rect -4886 617576 588810 617758
rect -2966 614294 586890 614476
rect -2966 614058 -1974 614294
rect -1738 614058 -1654 614294
rect -1418 614058 986 614294
rect 1222 614058 36986 614294
rect 37222 614058 72986 614294
rect 73222 614058 108986 614294
rect 109222 614058 144986 614294
rect 145222 614058 180986 614294
rect 181222 614058 216986 614294
rect 217222 614058 252986 614294
rect 253222 614058 288986 614294
rect 289222 614058 324986 614294
rect 325222 614058 360986 614294
rect 361222 614058 396986 614294
rect 397222 614058 432986 614294
rect 433222 614058 468986 614294
rect 469222 614058 504986 614294
rect 505222 614058 540986 614294
rect 541222 614058 576986 614294
rect 577222 614058 585342 614294
rect 585578 614058 585662 614294
rect 585898 614058 586890 614294
rect -2966 613876 586890 614058
rect -8726 607394 592650 607576
rect -8726 607158 -8694 607394
rect -8458 607158 -8374 607394
rect -8138 607158 30086 607394
rect 30322 607158 66086 607394
rect 66322 607158 102086 607394
rect 102322 607158 138086 607394
rect 138322 607158 174086 607394
rect 174322 607158 210086 607394
rect 210322 607158 246086 607394
rect 246322 607158 282086 607394
rect 282322 607158 318086 607394
rect 318322 607158 354086 607394
rect 354322 607158 390086 607394
rect 390322 607158 426086 607394
rect 426322 607158 462086 607394
rect 462322 607158 498086 607394
rect 498322 607158 534086 607394
rect 534322 607158 570086 607394
rect 570322 607158 592062 607394
rect 592298 607158 592382 607394
rect 592618 607158 592650 607394
rect -8726 606976 592650 607158
rect -6806 603694 590730 603876
rect -6806 603458 -6774 603694
rect -6538 603458 -6454 603694
rect -6218 603458 26386 603694
rect 26622 603458 62386 603694
rect 62622 603458 98386 603694
rect 98622 603458 134386 603694
rect 134622 603458 170386 603694
rect 170622 603458 206386 603694
rect 206622 603458 242386 603694
rect 242622 603458 278386 603694
rect 278622 603458 314386 603694
rect 314622 603458 350386 603694
rect 350622 603458 386386 603694
rect 386622 603458 422386 603694
rect 422622 603458 458386 603694
rect 458622 603458 494386 603694
rect 494622 603458 530386 603694
rect 530622 603458 566386 603694
rect 566622 603458 590142 603694
rect 590378 603458 590462 603694
rect 590698 603458 590730 603694
rect -6806 603276 590730 603458
rect -4886 599994 588810 600176
rect -4886 599758 -4854 599994
rect -4618 599758 -4534 599994
rect -4298 599758 22686 599994
rect 22922 599758 58686 599994
rect 58922 599758 94686 599994
rect 94922 599758 130686 599994
rect 130922 599758 166686 599994
rect 166922 599758 202686 599994
rect 202922 599758 238686 599994
rect 238922 599758 274686 599994
rect 274922 599758 310686 599994
rect 310922 599758 346686 599994
rect 346922 599758 382686 599994
rect 382922 599758 418686 599994
rect 418922 599758 454686 599994
rect 454922 599758 490686 599994
rect 490922 599758 526686 599994
rect 526922 599758 562686 599994
rect 562922 599758 588222 599994
rect 588458 599758 588542 599994
rect 588778 599758 588810 599994
rect -4886 599576 588810 599758
rect -2966 596294 586890 596476
rect -2966 596058 -2934 596294
rect -2698 596058 -2614 596294
rect -2378 596058 18986 596294
rect 19222 596058 54986 596294
rect 55222 596058 90986 596294
rect 91222 596058 126986 596294
rect 127222 596058 162986 596294
rect 163222 596058 198986 596294
rect 199222 596058 234986 596294
rect 235222 596058 270986 596294
rect 271222 596058 306986 596294
rect 307222 596058 342986 596294
rect 343222 596058 378986 596294
rect 379222 596058 414986 596294
rect 415222 596058 450986 596294
rect 451222 596058 486986 596294
rect 487222 596058 522986 596294
rect 523222 596058 558986 596294
rect 559222 596058 586302 596294
rect 586538 596058 586622 596294
rect 586858 596058 586890 596294
rect -2966 595876 586890 596058
rect -8726 589394 592650 589576
rect -8726 589158 -7734 589394
rect -7498 589158 -7414 589394
rect -7178 589158 12086 589394
rect 12322 589158 48086 589394
rect 48322 589158 84086 589394
rect 84322 589158 120086 589394
rect 120322 589158 156086 589394
rect 156322 589158 192086 589394
rect 192322 589158 228086 589394
rect 228322 589158 264086 589394
rect 264322 589158 300086 589394
rect 300322 589158 336086 589394
rect 336322 589158 372086 589394
rect 372322 589158 408086 589394
rect 408322 589158 444086 589394
rect 444322 589158 480086 589394
rect 480322 589158 516086 589394
rect 516322 589158 552086 589394
rect 552322 589158 591102 589394
rect 591338 589158 591422 589394
rect 591658 589158 592650 589394
rect -8726 588976 592650 589158
rect -6806 585694 590730 585876
rect -6806 585458 -5814 585694
rect -5578 585458 -5494 585694
rect -5258 585458 8386 585694
rect 8622 585458 44386 585694
rect 44622 585458 80386 585694
rect 80622 585458 116386 585694
rect 116622 585458 152386 585694
rect 152622 585458 188386 585694
rect 188622 585458 224386 585694
rect 224622 585458 260386 585694
rect 260622 585458 296386 585694
rect 296622 585458 332386 585694
rect 332622 585458 368386 585694
rect 368622 585458 404386 585694
rect 404622 585458 440386 585694
rect 440622 585458 476386 585694
rect 476622 585458 512386 585694
rect 512622 585458 548386 585694
rect 548622 585458 589182 585694
rect 589418 585458 589502 585694
rect 589738 585458 590730 585694
rect -6806 585276 590730 585458
rect -4886 581994 588810 582176
rect -4886 581758 -3894 581994
rect -3658 581758 -3574 581994
rect -3338 581758 4686 581994
rect 4922 581758 40686 581994
rect 40922 581758 76686 581994
rect 76922 581758 112686 581994
rect 112922 581758 148686 581994
rect 148922 581758 184686 581994
rect 184922 581758 220686 581994
rect 220922 581758 256686 581994
rect 256922 581758 292686 581994
rect 292922 581758 328686 581994
rect 328922 581758 364686 581994
rect 364922 581758 400686 581994
rect 400922 581758 436686 581994
rect 436922 581758 472686 581994
rect 472922 581758 508686 581994
rect 508922 581758 544686 581994
rect 544922 581758 580686 581994
rect 580922 581758 587262 581994
rect 587498 581758 587582 581994
rect 587818 581758 588810 581994
rect -4886 581576 588810 581758
rect -2966 578294 586890 578476
rect -2966 578058 -1974 578294
rect -1738 578058 -1654 578294
rect -1418 578058 986 578294
rect 1222 578058 36986 578294
rect 37222 578058 72986 578294
rect 73222 578058 108986 578294
rect 109222 578058 144986 578294
rect 145222 578058 180986 578294
rect 181222 578058 216986 578294
rect 217222 578058 252986 578294
rect 253222 578058 288986 578294
rect 289222 578058 324986 578294
rect 325222 578058 360986 578294
rect 361222 578058 396986 578294
rect 397222 578058 432986 578294
rect 433222 578058 468986 578294
rect 469222 578058 504986 578294
rect 505222 578058 540986 578294
rect 541222 578058 576986 578294
rect 577222 578058 585342 578294
rect 585578 578058 585662 578294
rect 585898 578058 586890 578294
rect -2966 577876 586890 578058
rect -8726 571394 592650 571576
rect -8726 571158 -8694 571394
rect -8458 571158 -8374 571394
rect -8138 571158 30086 571394
rect 30322 571158 66086 571394
rect 66322 571158 102086 571394
rect 102322 571158 138086 571394
rect 138322 571158 174086 571394
rect 174322 571158 210086 571394
rect 210322 571158 246086 571394
rect 246322 571158 282086 571394
rect 282322 571158 318086 571394
rect 318322 571158 354086 571394
rect 354322 571158 390086 571394
rect 390322 571158 426086 571394
rect 426322 571158 462086 571394
rect 462322 571158 498086 571394
rect 498322 571158 534086 571394
rect 534322 571158 570086 571394
rect 570322 571158 592062 571394
rect 592298 571158 592382 571394
rect 592618 571158 592650 571394
rect -8726 570976 592650 571158
rect -6806 567694 590730 567876
rect -6806 567458 -6774 567694
rect -6538 567458 -6454 567694
rect -6218 567458 26386 567694
rect 26622 567458 62386 567694
rect 62622 567458 98386 567694
rect 98622 567458 134386 567694
rect 134622 567458 170386 567694
rect 170622 567458 206386 567694
rect 206622 567458 242386 567694
rect 242622 567458 278386 567694
rect 278622 567458 314386 567694
rect 314622 567458 350386 567694
rect 350622 567458 386386 567694
rect 386622 567458 422386 567694
rect 422622 567458 458386 567694
rect 458622 567458 494386 567694
rect 494622 567458 530386 567694
rect 530622 567458 566386 567694
rect 566622 567458 590142 567694
rect 590378 567458 590462 567694
rect 590698 567458 590730 567694
rect -6806 567276 590730 567458
rect -4886 563994 588810 564176
rect -4886 563758 -4854 563994
rect -4618 563758 -4534 563994
rect -4298 563758 22686 563994
rect 22922 563758 58686 563994
rect 58922 563758 94686 563994
rect 94922 563758 130686 563994
rect 130922 563758 166686 563994
rect 166922 563758 202686 563994
rect 202922 563758 238686 563994
rect 238922 563758 274686 563994
rect 274922 563758 310686 563994
rect 310922 563758 346686 563994
rect 346922 563758 382686 563994
rect 382922 563758 418686 563994
rect 418922 563758 454686 563994
rect 454922 563758 490686 563994
rect 490922 563758 526686 563994
rect 526922 563758 562686 563994
rect 562922 563758 588222 563994
rect 588458 563758 588542 563994
rect 588778 563758 588810 563994
rect -4886 563576 588810 563758
rect -2966 560294 586890 560476
rect -2966 560058 -2934 560294
rect -2698 560058 -2614 560294
rect -2378 560058 18986 560294
rect 19222 560058 54986 560294
rect 55222 560058 90986 560294
rect 91222 560058 126986 560294
rect 127222 560058 162986 560294
rect 163222 560058 198986 560294
rect 199222 560058 234986 560294
rect 235222 560058 270986 560294
rect 271222 560058 306986 560294
rect 307222 560058 342986 560294
rect 343222 560058 378986 560294
rect 379222 560058 414986 560294
rect 415222 560058 450986 560294
rect 451222 560058 486986 560294
rect 487222 560058 522986 560294
rect 523222 560058 558986 560294
rect 559222 560058 586302 560294
rect 586538 560058 586622 560294
rect 586858 560058 586890 560294
rect -2966 559876 586890 560058
rect -8726 553394 592650 553576
rect -8726 553158 -7734 553394
rect -7498 553158 -7414 553394
rect -7178 553158 12086 553394
rect 12322 553158 48086 553394
rect 48322 553158 84086 553394
rect 84322 553158 120086 553394
rect 120322 553158 156086 553394
rect 156322 553158 192086 553394
rect 192322 553158 228086 553394
rect 228322 553158 264086 553394
rect 264322 553158 300086 553394
rect 300322 553158 336086 553394
rect 336322 553158 372086 553394
rect 372322 553158 408086 553394
rect 408322 553158 444086 553394
rect 444322 553158 480086 553394
rect 480322 553158 516086 553394
rect 516322 553158 552086 553394
rect 552322 553158 591102 553394
rect 591338 553158 591422 553394
rect 591658 553158 592650 553394
rect -8726 552976 592650 553158
rect -6806 549694 590730 549876
rect -6806 549458 -5814 549694
rect -5578 549458 -5494 549694
rect -5258 549458 8386 549694
rect 8622 549458 44386 549694
rect 44622 549458 80386 549694
rect 80622 549458 116386 549694
rect 116622 549458 152386 549694
rect 152622 549458 188386 549694
rect 188622 549458 224386 549694
rect 224622 549458 260386 549694
rect 260622 549458 296386 549694
rect 296622 549458 332386 549694
rect 332622 549458 368386 549694
rect 368622 549458 404386 549694
rect 404622 549458 440386 549694
rect 440622 549458 476386 549694
rect 476622 549458 512386 549694
rect 512622 549458 548386 549694
rect 548622 549458 589182 549694
rect 589418 549458 589502 549694
rect 589738 549458 590730 549694
rect -6806 549276 590730 549458
rect -4886 545994 588810 546176
rect -4886 545758 -3894 545994
rect -3658 545758 -3574 545994
rect -3338 545758 4686 545994
rect 4922 545758 40686 545994
rect 40922 545758 76686 545994
rect 76922 545758 112686 545994
rect 112922 545758 148686 545994
rect 148922 545758 184686 545994
rect 184922 545758 220686 545994
rect 220922 545758 256686 545994
rect 256922 545758 292686 545994
rect 292922 545758 328686 545994
rect 328922 545758 364686 545994
rect 364922 545758 400686 545994
rect 400922 545758 436686 545994
rect 436922 545758 472686 545994
rect 472922 545758 508686 545994
rect 508922 545758 544686 545994
rect 544922 545758 580686 545994
rect 580922 545758 587262 545994
rect 587498 545758 587582 545994
rect 587818 545758 588810 545994
rect -4886 545576 588810 545758
rect -2966 542294 586890 542476
rect -2966 542058 -1974 542294
rect -1738 542058 -1654 542294
rect -1418 542058 986 542294
rect 1222 542058 36986 542294
rect 37222 542058 72986 542294
rect 73222 542058 108986 542294
rect 109222 542058 144986 542294
rect 145222 542058 180986 542294
rect 181222 542058 216986 542294
rect 217222 542058 252986 542294
rect 253222 542058 288986 542294
rect 289222 542058 324986 542294
rect 325222 542058 360986 542294
rect 361222 542058 396986 542294
rect 397222 542058 432986 542294
rect 433222 542058 468986 542294
rect 469222 542058 504986 542294
rect 505222 542058 540986 542294
rect 541222 542058 576986 542294
rect 577222 542058 585342 542294
rect 585578 542058 585662 542294
rect 585898 542058 586890 542294
rect -2966 541876 586890 542058
rect -8726 535394 592650 535576
rect -8726 535158 -8694 535394
rect -8458 535158 -8374 535394
rect -8138 535158 30086 535394
rect 30322 535158 66086 535394
rect 66322 535158 102086 535394
rect 102322 535158 138086 535394
rect 138322 535158 174086 535394
rect 174322 535158 210086 535394
rect 210322 535158 246086 535394
rect 246322 535158 282086 535394
rect 282322 535158 318086 535394
rect 318322 535158 354086 535394
rect 354322 535158 390086 535394
rect 390322 535158 426086 535394
rect 426322 535158 462086 535394
rect 462322 535158 498086 535394
rect 498322 535158 534086 535394
rect 534322 535158 570086 535394
rect 570322 535158 592062 535394
rect 592298 535158 592382 535394
rect 592618 535158 592650 535394
rect -8726 534976 592650 535158
rect -6806 531694 590730 531876
rect -6806 531458 -6774 531694
rect -6538 531458 -6454 531694
rect -6218 531458 26386 531694
rect 26622 531458 62386 531694
rect 62622 531458 98386 531694
rect 98622 531458 134386 531694
rect 134622 531458 170386 531694
rect 170622 531458 206386 531694
rect 206622 531458 242386 531694
rect 242622 531458 278386 531694
rect 278622 531458 314386 531694
rect 314622 531458 350386 531694
rect 350622 531458 386386 531694
rect 386622 531458 422386 531694
rect 422622 531458 458386 531694
rect 458622 531458 494386 531694
rect 494622 531458 530386 531694
rect 530622 531458 566386 531694
rect 566622 531458 590142 531694
rect 590378 531458 590462 531694
rect 590698 531458 590730 531694
rect -6806 531276 590730 531458
rect -4886 527994 588810 528176
rect -4886 527758 -4854 527994
rect -4618 527758 -4534 527994
rect -4298 527758 22686 527994
rect 22922 527758 58686 527994
rect 58922 527758 94686 527994
rect 94922 527758 130686 527994
rect 130922 527758 166686 527994
rect 166922 527758 202686 527994
rect 202922 527758 238686 527994
rect 238922 527758 274686 527994
rect 274922 527758 310686 527994
rect 310922 527758 346686 527994
rect 346922 527758 382686 527994
rect 382922 527758 418686 527994
rect 418922 527758 454686 527994
rect 454922 527758 490686 527994
rect 490922 527758 526686 527994
rect 526922 527758 562686 527994
rect 562922 527758 588222 527994
rect 588458 527758 588542 527994
rect 588778 527758 588810 527994
rect -4886 527576 588810 527758
rect -2966 524294 586890 524476
rect -2966 524058 -2934 524294
rect -2698 524058 -2614 524294
rect -2378 524058 18986 524294
rect 19222 524058 54986 524294
rect 55222 524058 90986 524294
rect 91222 524058 126986 524294
rect 127222 524058 162986 524294
rect 163222 524058 198986 524294
rect 199222 524058 234986 524294
rect 235222 524058 270986 524294
rect 271222 524058 306986 524294
rect 307222 524058 342986 524294
rect 343222 524058 378986 524294
rect 379222 524058 414986 524294
rect 415222 524058 450986 524294
rect 451222 524058 486986 524294
rect 487222 524058 522986 524294
rect 523222 524058 558986 524294
rect 559222 524058 586302 524294
rect 586538 524058 586622 524294
rect 586858 524058 586890 524294
rect -2966 523876 586890 524058
rect -8726 517394 592650 517576
rect -8726 517158 -7734 517394
rect -7498 517158 -7414 517394
rect -7178 517158 12086 517394
rect 12322 517158 48086 517394
rect 48322 517158 84086 517394
rect 84322 517158 120086 517394
rect 120322 517158 156086 517394
rect 156322 517158 192086 517394
rect 192322 517158 228086 517394
rect 228322 517158 264086 517394
rect 264322 517158 300086 517394
rect 300322 517158 336086 517394
rect 336322 517158 372086 517394
rect 372322 517158 408086 517394
rect 408322 517158 444086 517394
rect 444322 517158 480086 517394
rect 480322 517158 516086 517394
rect 516322 517158 552086 517394
rect 552322 517158 591102 517394
rect 591338 517158 591422 517394
rect 591658 517158 592650 517394
rect -8726 516976 592650 517158
rect -6806 513694 590730 513876
rect -6806 513458 -5814 513694
rect -5578 513458 -5494 513694
rect -5258 513458 8386 513694
rect 8622 513458 44386 513694
rect 44622 513458 80386 513694
rect 80622 513458 116386 513694
rect 116622 513458 152386 513694
rect 152622 513458 188386 513694
rect 188622 513458 224386 513694
rect 224622 513458 260386 513694
rect 260622 513458 296386 513694
rect 296622 513458 332386 513694
rect 332622 513458 368386 513694
rect 368622 513458 404386 513694
rect 404622 513458 440386 513694
rect 440622 513458 476386 513694
rect 476622 513458 512386 513694
rect 512622 513458 548386 513694
rect 548622 513458 589182 513694
rect 589418 513458 589502 513694
rect 589738 513458 590730 513694
rect -6806 513276 590730 513458
rect -4886 509994 588810 510176
rect -4886 509758 -3894 509994
rect -3658 509758 -3574 509994
rect -3338 509758 4686 509994
rect 4922 509758 40686 509994
rect 40922 509758 76686 509994
rect 76922 509758 112686 509994
rect 112922 509758 148686 509994
rect 148922 509758 184686 509994
rect 184922 509758 220686 509994
rect 220922 509758 256686 509994
rect 256922 509758 292686 509994
rect 292922 509758 328686 509994
rect 328922 509758 364686 509994
rect 364922 509758 400686 509994
rect 400922 509758 436686 509994
rect 436922 509758 472686 509994
rect 472922 509758 508686 509994
rect 508922 509758 544686 509994
rect 544922 509758 580686 509994
rect 580922 509758 587262 509994
rect 587498 509758 587582 509994
rect 587818 509758 588810 509994
rect -4886 509576 588810 509758
rect -2966 506294 586890 506476
rect -2966 506058 -1974 506294
rect -1738 506058 -1654 506294
rect -1418 506058 986 506294
rect 1222 506058 36986 506294
rect 37222 506058 72986 506294
rect 73222 506058 108986 506294
rect 109222 506058 144986 506294
rect 145222 506058 180986 506294
rect 181222 506058 216986 506294
rect 217222 506058 252986 506294
rect 253222 506058 288986 506294
rect 289222 506058 324986 506294
rect 325222 506058 360986 506294
rect 361222 506058 396986 506294
rect 397222 506058 432986 506294
rect 433222 506058 468986 506294
rect 469222 506058 504986 506294
rect 505222 506058 540986 506294
rect 541222 506058 576986 506294
rect 577222 506058 585342 506294
rect 585578 506058 585662 506294
rect 585898 506058 586890 506294
rect -2966 505876 586890 506058
rect -8726 499394 592650 499576
rect -8726 499158 -8694 499394
rect -8458 499158 -8374 499394
rect -8138 499158 30086 499394
rect 30322 499158 66086 499394
rect 66322 499158 102086 499394
rect 102322 499158 138086 499394
rect 138322 499158 174086 499394
rect 174322 499158 210086 499394
rect 210322 499158 246086 499394
rect 246322 499158 282086 499394
rect 282322 499158 318086 499394
rect 318322 499158 354086 499394
rect 354322 499158 390086 499394
rect 390322 499158 426086 499394
rect 426322 499158 462086 499394
rect 462322 499158 498086 499394
rect 498322 499158 534086 499394
rect 534322 499158 570086 499394
rect 570322 499158 592062 499394
rect 592298 499158 592382 499394
rect 592618 499158 592650 499394
rect -8726 498976 592650 499158
rect -6806 495694 590730 495876
rect -6806 495458 -6774 495694
rect -6538 495458 -6454 495694
rect -6218 495458 26386 495694
rect 26622 495458 62386 495694
rect 62622 495458 98386 495694
rect 98622 495458 134386 495694
rect 134622 495458 170386 495694
rect 170622 495458 206386 495694
rect 206622 495458 242386 495694
rect 242622 495458 278386 495694
rect 278622 495458 314386 495694
rect 314622 495458 350386 495694
rect 350622 495458 386386 495694
rect 386622 495458 422386 495694
rect 422622 495458 458386 495694
rect 458622 495458 494386 495694
rect 494622 495458 530386 495694
rect 530622 495458 566386 495694
rect 566622 495458 590142 495694
rect 590378 495458 590462 495694
rect 590698 495458 590730 495694
rect -6806 495276 590730 495458
rect -4886 491994 588810 492176
rect -4886 491758 -4854 491994
rect -4618 491758 -4534 491994
rect -4298 491758 22686 491994
rect 22922 491758 58686 491994
rect 58922 491758 94686 491994
rect 94922 491758 130686 491994
rect 130922 491758 166686 491994
rect 166922 491758 202686 491994
rect 202922 491758 238686 491994
rect 238922 491758 274686 491994
rect 274922 491758 310686 491994
rect 310922 491758 346686 491994
rect 346922 491758 382686 491994
rect 382922 491758 418686 491994
rect 418922 491758 454686 491994
rect 454922 491758 490686 491994
rect 490922 491758 526686 491994
rect 526922 491758 562686 491994
rect 562922 491758 588222 491994
rect 588458 491758 588542 491994
rect 588778 491758 588810 491994
rect -4886 491576 588810 491758
rect -2966 488294 586890 488476
rect -2966 488058 -2934 488294
rect -2698 488058 -2614 488294
rect -2378 488058 18986 488294
rect 19222 488058 54986 488294
rect 55222 488058 90986 488294
rect 91222 488058 126986 488294
rect 127222 488058 162986 488294
rect 163222 488058 198986 488294
rect 199222 488058 234986 488294
rect 235222 488058 270986 488294
rect 271222 488058 306986 488294
rect 307222 488058 342986 488294
rect 343222 488058 378986 488294
rect 379222 488058 414986 488294
rect 415222 488058 450986 488294
rect 451222 488058 486986 488294
rect 487222 488058 522986 488294
rect 523222 488058 558986 488294
rect 559222 488058 586302 488294
rect 586538 488058 586622 488294
rect 586858 488058 586890 488294
rect -2966 487876 586890 488058
rect -8726 481394 592650 481576
rect -8726 481158 -7734 481394
rect -7498 481158 -7414 481394
rect -7178 481158 12086 481394
rect 12322 481158 48086 481394
rect 48322 481158 84086 481394
rect 84322 481158 120086 481394
rect 120322 481158 156086 481394
rect 156322 481158 192086 481394
rect 192322 481158 228086 481394
rect 228322 481158 264086 481394
rect 264322 481158 300086 481394
rect 300322 481158 336086 481394
rect 336322 481158 372086 481394
rect 372322 481158 408086 481394
rect 408322 481158 444086 481394
rect 444322 481158 480086 481394
rect 480322 481158 516086 481394
rect 516322 481158 552086 481394
rect 552322 481158 591102 481394
rect 591338 481158 591422 481394
rect 591658 481158 592650 481394
rect -8726 480976 592650 481158
rect -6806 477694 590730 477876
rect -6806 477458 -5814 477694
rect -5578 477458 -5494 477694
rect -5258 477458 8386 477694
rect 8622 477458 44386 477694
rect 44622 477458 80386 477694
rect 80622 477458 116386 477694
rect 116622 477458 152386 477694
rect 152622 477458 188386 477694
rect 188622 477458 224386 477694
rect 224622 477458 260386 477694
rect 260622 477458 296386 477694
rect 296622 477458 332386 477694
rect 332622 477458 368386 477694
rect 368622 477458 404386 477694
rect 404622 477458 440386 477694
rect 440622 477458 476386 477694
rect 476622 477458 512386 477694
rect 512622 477458 548386 477694
rect 548622 477458 589182 477694
rect 589418 477458 589502 477694
rect 589738 477458 590730 477694
rect -6806 477276 590730 477458
rect -4886 473994 588810 474176
rect -4886 473758 -3894 473994
rect -3658 473758 -3574 473994
rect -3338 473758 4686 473994
rect 4922 473758 40686 473994
rect 40922 473758 76686 473994
rect 76922 473758 112686 473994
rect 112922 473758 148686 473994
rect 148922 473758 184686 473994
rect 184922 473758 220686 473994
rect 220922 473758 256686 473994
rect 256922 473758 292686 473994
rect 292922 473758 328686 473994
rect 328922 473758 364686 473994
rect 364922 473758 400686 473994
rect 400922 473758 436686 473994
rect 436922 473758 472686 473994
rect 472922 473758 508686 473994
rect 508922 473758 544686 473994
rect 544922 473758 580686 473994
rect 580922 473758 587262 473994
rect 587498 473758 587582 473994
rect 587818 473758 588810 473994
rect -4886 473576 588810 473758
rect -2966 470294 586890 470476
rect -2966 470058 -1974 470294
rect -1738 470058 -1654 470294
rect -1418 470058 986 470294
rect 1222 470058 36986 470294
rect 37222 470058 72986 470294
rect 73222 470058 108986 470294
rect 109222 470058 144986 470294
rect 145222 470058 180986 470294
rect 181222 470058 216986 470294
rect 217222 470058 252986 470294
rect 253222 470058 288986 470294
rect 289222 470058 324986 470294
rect 325222 470058 360986 470294
rect 361222 470058 396986 470294
rect 397222 470058 432986 470294
rect 433222 470058 468986 470294
rect 469222 470058 504986 470294
rect 505222 470058 540986 470294
rect 541222 470058 576986 470294
rect 577222 470058 585342 470294
rect 585578 470058 585662 470294
rect 585898 470058 586890 470294
rect -2966 469876 586890 470058
rect -8726 463394 592650 463576
rect -8726 463158 -8694 463394
rect -8458 463158 -8374 463394
rect -8138 463158 30086 463394
rect 30322 463158 66086 463394
rect 66322 463158 102086 463394
rect 102322 463158 138086 463394
rect 138322 463158 174086 463394
rect 174322 463158 210086 463394
rect 210322 463158 246086 463394
rect 246322 463158 282086 463394
rect 282322 463158 318086 463394
rect 318322 463158 354086 463394
rect 354322 463158 390086 463394
rect 390322 463158 426086 463394
rect 426322 463158 462086 463394
rect 462322 463158 498086 463394
rect 498322 463158 534086 463394
rect 534322 463158 570086 463394
rect 570322 463158 592062 463394
rect 592298 463158 592382 463394
rect 592618 463158 592650 463394
rect -8726 462976 592650 463158
rect -6806 459694 590730 459876
rect -6806 459458 -6774 459694
rect -6538 459458 -6454 459694
rect -6218 459458 26386 459694
rect 26622 459458 62386 459694
rect 62622 459458 98386 459694
rect 98622 459458 134386 459694
rect 134622 459458 170386 459694
rect 170622 459458 206386 459694
rect 206622 459458 242386 459694
rect 242622 459458 278386 459694
rect 278622 459458 314386 459694
rect 314622 459458 350386 459694
rect 350622 459458 386386 459694
rect 386622 459458 422386 459694
rect 422622 459458 458386 459694
rect 458622 459458 494386 459694
rect 494622 459458 530386 459694
rect 530622 459458 566386 459694
rect 566622 459458 590142 459694
rect 590378 459458 590462 459694
rect 590698 459458 590730 459694
rect -6806 459276 590730 459458
rect -4886 455994 588810 456176
rect -4886 455758 -4854 455994
rect -4618 455758 -4534 455994
rect -4298 455758 22686 455994
rect 22922 455758 58686 455994
rect 58922 455758 94686 455994
rect 94922 455758 130686 455994
rect 130922 455758 166686 455994
rect 166922 455758 202686 455994
rect 202922 455758 238686 455994
rect 238922 455758 274686 455994
rect 274922 455758 310686 455994
rect 310922 455758 346686 455994
rect 346922 455758 382686 455994
rect 382922 455758 418686 455994
rect 418922 455758 454686 455994
rect 454922 455758 490686 455994
rect 490922 455758 526686 455994
rect 526922 455758 562686 455994
rect 562922 455758 588222 455994
rect 588458 455758 588542 455994
rect 588778 455758 588810 455994
rect -4886 455576 588810 455758
rect -2966 452294 586890 452476
rect -2966 452058 -2934 452294
rect -2698 452058 -2614 452294
rect -2378 452058 18986 452294
rect 19222 452058 54986 452294
rect 55222 452058 90986 452294
rect 91222 452058 126986 452294
rect 127222 452058 162986 452294
rect 163222 452058 198986 452294
rect 199222 452058 234986 452294
rect 235222 452058 270986 452294
rect 271222 452058 306986 452294
rect 307222 452058 342986 452294
rect 343222 452058 378986 452294
rect 379222 452058 414986 452294
rect 415222 452058 450986 452294
rect 451222 452058 486986 452294
rect 487222 452058 522986 452294
rect 523222 452058 558986 452294
rect 559222 452058 586302 452294
rect 586538 452058 586622 452294
rect 586858 452058 586890 452294
rect -2966 451876 586890 452058
rect -8726 445394 592650 445576
rect -8726 445158 -7734 445394
rect -7498 445158 -7414 445394
rect -7178 445158 12086 445394
rect 12322 445158 48086 445394
rect 48322 445158 84086 445394
rect 84322 445158 120086 445394
rect 120322 445158 156086 445394
rect 156322 445158 192086 445394
rect 192322 445158 228086 445394
rect 228322 445158 264086 445394
rect 264322 445158 300086 445394
rect 300322 445158 336086 445394
rect 336322 445158 372086 445394
rect 372322 445158 408086 445394
rect 408322 445158 444086 445394
rect 444322 445158 480086 445394
rect 480322 445158 516086 445394
rect 516322 445158 552086 445394
rect 552322 445158 591102 445394
rect 591338 445158 591422 445394
rect 591658 445158 592650 445394
rect -8726 444976 592650 445158
rect -6806 441694 590730 441876
rect -6806 441458 -5814 441694
rect -5578 441458 -5494 441694
rect -5258 441458 8386 441694
rect 8622 441458 44386 441694
rect 44622 441458 80386 441694
rect 80622 441458 116386 441694
rect 116622 441458 152386 441694
rect 152622 441458 188386 441694
rect 188622 441458 224386 441694
rect 224622 441458 260386 441694
rect 260622 441458 296386 441694
rect 296622 441458 332386 441694
rect 332622 441458 368386 441694
rect 368622 441458 404386 441694
rect 404622 441458 440386 441694
rect 440622 441458 476386 441694
rect 476622 441458 512386 441694
rect 512622 441458 548386 441694
rect 548622 441458 589182 441694
rect 589418 441458 589502 441694
rect 589738 441458 590730 441694
rect -6806 441276 590730 441458
rect -4886 437994 588810 438176
rect -4886 437758 -3894 437994
rect -3658 437758 -3574 437994
rect -3338 437758 4686 437994
rect 4922 437758 40686 437994
rect 40922 437758 76686 437994
rect 76922 437758 112686 437994
rect 112922 437758 148686 437994
rect 148922 437758 184686 437994
rect 184922 437758 220686 437994
rect 220922 437758 256686 437994
rect 256922 437758 292686 437994
rect 292922 437758 328686 437994
rect 328922 437758 364686 437994
rect 364922 437758 400686 437994
rect 400922 437758 436686 437994
rect 436922 437758 472686 437994
rect 472922 437758 508686 437994
rect 508922 437758 544686 437994
rect 544922 437758 580686 437994
rect 580922 437758 587262 437994
rect 587498 437758 587582 437994
rect 587818 437758 588810 437994
rect -4886 437576 588810 437758
rect -2966 434294 586890 434476
rect -2966 434058 -1974 434294
rect -1738 434058 -1654 434294
rect -1418 434058 986 434294
rect 1222 434058 36986 434294
rect 37222 434058 72986 434294
rect 73222 434058 108986 434294
rect 109222 434058 144986 434294
rect 145222 434058 180986 434294
rect 181222 434058 216986 434294
rect 217222 434058 252986 434294
rect 253222 434058 288986 434294
rect 289222 434058 324986 434294
rect 325222 434058 360986 434294
rect 361222 434058 396986 434294
rect 397222 434058 432986 434294
rect 433222 434058 468986 434294
rect 469222 434058 504986 434294
rect 505222 434058 540986 434294
rect 541222 434058 576986 434294
rect 577222 434058 585342 434294
rect 585578 434058 585662 434294
rect 585898 434058 586890 434294
rect -2966 433876 586890 434058
rect -8726 427394 592650 427576
rect -8726 427158 -8694 427394
rect -8458 427158 -8374 427394
rect -8138 427158 30086 427394
rect 30322 427158 66086 427394
rect 66322 427158 102086 427394
rect 102322 427158 138086 427394
rect 138322 427158 174086 427394
rect 174322 427158 210086 427394
rect 210322 427158 246086 427394
rect 246322 427158 282086 427394
rect 282322 427158 318086 427394
rect 318322 427158 354086 427394
rect 354322 427158 390086 427394
rect 390322 427158 426086 427394
rect 426322 427158 462086 427394
rect 462322 427158 498086 427394
rect 498322 427158 534086 427394
rect 534322 427158 570086 427394
rect 570322 427158 592062 427394
rect 592298 427158 592382 427394
rect 592618 427158 592650 427394
rect -8726 426976 592650 427158
rect -6806 423694 590730 423876
rect -6806 423458 -6774 423694
rect -6538 423458 -6454 423694
rect -6218 423458 26386 423694
rect 26622 423458 206386 423694
rect 206622 423458 242386 423694
rect 242622 423458 278386 423694
rect 278622 423458 314386 423694
rect 314622 423458 494386 423694
rect 494622 423458 530386 423694
rect 530622 423458 566386 423694
rect 566622 423458 590142 423694
rect 590378 423458 590462 423694
rect 590698 423458 590730 423694
rect -6806 423276 590730 423458
rect -4886 419994 588810 420176
rect -4886 419758 -4854 419994
rect -4618 419758 -4534 419994
rect -4298 419758 22686 419994
rect 22922 419758 202686 419994
rect 202922 419758 238686 419994
rect 238922 419758 274686 419994
rect 274922 419758 310686 419994
rect 310922 419758 490686 419994
rect 490922 419758 526686 419994
rect 526922 419758 562686 419994
rect 562922 419758 588222 419994
rect 588458 419758 588542 419994
rect 588778 419758 588810 419994
rect -4886 419576 588810 419758
rect -2966 416294 586890 416476
rect -2966 416058 -2934 416294
rect -2698 416058 -2614 416294
rect -2378 416058 18986 416294
rect 19222 416058 40328 416294
rect 40564 416058 176056 416294
rect 176292 416058 198986 416294
rect 199222 416058 234986 416294
rect 235222 416058 270986 416294
rect 271222 416058 306986 416294
rect 307222 416058 340328 416294
rect 340564 416058 476056 416294
rect 476292 416058 486986 416294
rect 487222 416058 522986 416294
rect 523222 416058 558986 416294
rect 559222 416058 586302 416294
rect 586538 416058 586622 416294
rect 586858 416058 586890 416294
rect -2966 415876 586890 416058
rect -8726 409394 592650 409576
rect -8726 409158 -7734 409394
rect -7498 409158 -7414 409394
rect -7178 409158 12086 409394
rect 12322 409158 192086 409394
rect 192322 409158 228086 409394
rect 228322 409158 264086 409394
rect 264322 409158 300086 409394
rect 300322 409158 336086 409394
rect 336322 409158 480086 409394
rect 480322 409158 516086 409394
rect 516322 409158 552086 409394
rect 552322 409158 591102 409394
rect 591338 409158 591422 409394
rect 591658 409158 592650 409394
rect -8726 408976 592650 409158
rect -6806 405694 590730 405876
rect -6806 405458 -5814 405694
rect -5578 405458 -5494 405694
rect -5258 405458 8386 405694
rect 8622 405458 188386 405694
rect 188622 405458 224386 405694
rect 224622 405458 260386 405694
rect 260622 405458 296386 405694
rect 296622 405458 332386 405694
rect 332622 405458 512386 405694
rect 512622 405458 548386 405694
rect 548622 405458 589182 405694
rect 589418 405458 589502 405694
rect 589738 405458 590730 405694
rect -6806 405276 590730 405458
rect -4886 401994 588810 402176
rect -4886 401758 -3894 401994
rect -3658 401758 -3574 401994
rect -3338 401758 4686 401994
rect 4922 401758 184686 401994
rect 184922 401758 220686 401994
rect 220922 401758 256686 401994
rect 256922 401758 292686 401994
rect 292922 401758 328686 401994
rect 328922 401758 508686 401994
rect 508922 401758 544686 401994
rect 544922 401758 580686 401994
rect 580922 401758 587262 401994
rect 587498 401758 587582 401994
rect 587818 401758 588810 401994
rect -4886 401576 588810 401758
rect -2966 398294 586890 398476
rect -2966 398058 -1974 398294
rect -1738 398058 -1654 398294
rect -1418 398058 986 398294
rect 1222 398058 36986 398294
rect 37222 398058 41008 398294
rect 41244 398058 175376 398294
rect 175612 398058 180986 398294
rect 181222 398058 216986 398294
rect 217222 398058 252986 398294
rect 253222 398058 288986 398294
rect 289222 398058 324986 398294
rect 325222 398058 341008 398294
rect 341244 398058 475376 398294
rect 475612 398058 504986 398294
rect 505222 398058 540986 398294
rect 541222 398058 576986 398294
rect 577222 398058 585342 398294
rect 585578 398058 585662 398294
rect 585898 398058 586890 398294
rect -2966 397876 586890 398058
rect -8726 391394 592650 391576
rect -8726 391158 -8694 391394
rect -8458 391158 -8374 391394
rect -8138 391158 30086 391394
rect 30322 391158 210086 391394
rect 210322 391158 246086 391394
rect 246322 391158 282086 391394
rect 282322 391158 318086 391394
rect 318322 391158 498086 391394
rect 498322 391158 534086 391394
rect 534322 391158 570086 391394
rect 570322 391158 592062 391394
rect 592298 391158 592382 391394
rect 592618 391158 592650 391394
rect -8726 390976 592650 391158
rect -6806 387694 590730 387876
rect -6806 387458 -6774 387694
rect -6538 387458 -6454 387694
rect -6218 387458 26386 387694
rect 26622 387458 206386 387694
rect 206622 387458 242386 387694
rect 242622 387458 278386 387694
rect 278622 387458 314386 387694
rect 314622 387458 494386 387694
rect 494622 387458 530386 387694
rect 530622 387458 566386 387694
rect 566622 387458 590142 387694
rect 590378 387458 590462 387694
rect 590698 387458 590730 387694
rect -6806 387276 590730 387458
rect -4886 383994 588810 384176
rect -4886 383758 -4854 383994
rect -4618 383758 -4534 383994
rect -4298 383758 22686 383994
rect 22922 383758 202686 383994
rect 202922 383758 238686 383994
rect 238922 383758 274686 383994
rect 274922 383758 310686 383994
rect 310922 383758 490686 383994
rect 490922 383758 526686 383994
rect 526922 383758 562686 383994
rect 562922 383758 588222 383994
rect 588458 383758 588542 383994
rect 588778 383758 588810 383994
rect -4886 383576 588810 383758
rect -2966 380294 586890 380476
rect -2966 380058 -2934 380294
rect -2698 380058 -2614 380294
rect -2378 380058 18986 380294
rect 19222 380058 40328 380294
rect 40564 380058 176056 380294
rect 176292 380058 198986 380294
rect 199222 380058 234986 380294
rect 235222 380058 270986 380294
rect 271222 380058 306986 380294
rect 307222 380058 340328 380294
rect 340564 380058 476056 380294
rect 476292 380058 486986 380294
rect 487222 380058 522986 380294
rect 523222 380058 558986 380294
rect 559222 380058 586302 380294
rect 586538 380058 586622 380294
rect 586858 380058 586890 380294
rect -2966 379876 586890 380058
rect -8726 373394 592650 373576
rect -8726 373158 -7734 373394
rect -7498 373158 -7414 373394
rect -7178 373158 12086 373394
rect 12322 373158 192086 373394
rect 192322 373158 228086 373394
rect 228322 373158 264086 373394
rect 264322 373158 300086 373394
rect 300322 373158 336086 373394
rect 336322 373158 480086 373394
rect 480322 373158 516086 373394
rect 516322 373158 552086 373394
rect 552322 373158 591102 373394
rect 591338 373158 591422 373394
rect 591658 373158 592650 373394
rect -8726 372976 592650 373158
rect -6806 369694 590730 369876
rect -6806 369458 -5814 369694
rect -5578 369458 -5494 369694
rect -5258 369458 8386 369694
rect 8622 369458 188386 369694
rect 188622 369458 224386 369694
rect 224622 369458 260386 369694
rect 260622 369458 296386 369694
rect 296622 369458 332386 369694
rect 332622 369458 512386 369694
rect 512622 369458 548386 369694
rect 548622 369458 589182 369694
rect 589418 369458 589502 369694
rect 589738 369458 590730 369694
rect -6806 369276 590730 369458
rect -4886 365994 588810 366176
rect -4886 365758 -3894 365994
rect -3658 365758 -3574 365994
rect -3338 365758 4686 365994
rect 4922 365758 184686 365994
rect 184922 365758 220686 365994
rect 220922 365758 256686 365994
rect 256922 365758 292686 365994
rect 292922 365758 328686 365994
rect 328922 365758 508686 365994
rect 508922 365758 544686 365994
rect 544922 365758 580686 365994
rect 580922 365758 587262 365994
rect 587498 365758 587582 365994
rect 587818 365758 588810 365994
rect -4886 365576 588810 365758
rect -2966 362294 586890 362476
rect -2966 362058 -1974 362294
rect -1738 362058 -1654 362294
rect -1418 362058 986 362294
rect 1222 362058 36986 362294
rect 37222 362058 41008 362294
rect 41244 362058 175376 362294
rect 175612 362058 180986 362294
rect 181222 362058 216986 362294
rect 217222 362058 252986 362294
rect 253222 362058 288986 362294
rect 289222 362058 324986 362294
rect 325222 362058 341008 362294
rect 341244 362058 475376 362294
rect 475612 362058 504986 362294
rect 505222 362058 540986 362294
rect 541222 362058 576986 362294
rect 577222 362058 585342 362294
rect 585578 362058 585662 362294
rect 585898 362058 586890 362294
rect -2966 361876 586890 362058
rect -8726 355394 592650 355576
rect -8726 355158 -8694 355394
rect -8458 355158 -8374 355394
rect -8138 355158 30086 355394
rect 30322 355158 210086 355394
rect 210322 355158 246086 355394
rect 246322 355158 282086 355394
rect 282322 355158 318086 355394
rect 318322 355158 498086 355394
rect 498322 355158 534086 355394
rect 534322 355158 570086 355394
rect 570322 355158 592062 355394
rect 592298 355158 592382 355394
rect 592618 355158 592650 355394
rect -8726 354976 592650 355158
rect -6806 351694 590730 351876
rect -6806 351458 -6774 351694
rect -6538 351458 -6454 351694
rect -6218 351458 26386 351694
rect 26622 351458 206386 351694
rect 206622 351458 242386 351694
rect 242622 351458 278386 351694
rect 278622 351458 314386 351694
rect 314622 351458 494386 351694
rect 494622 351458 530386 351694
rect 530622 351458 566386 351694
rect 566622 351458 590142 351694
rect 590378 351458 590462 351694
rect 590698 351458 590730 351694
rect -6806 351276 590730 351458
rect -4886 347994 588810 348176
rect -4886 347758 -4854 347994
rect -4618 347758 -4534 347994
rect -4298 347758 22686 347994
rect 22922 347758 202686 347994
rect 202922 347758 238686 347994
rect 238922 347758 274686 347994
rect 274922 347758 310686 347994
rect 310922 347758 490686 347994
rect 490922 347758 526686 347994
rect 526922 347758 562686 347994
rect 562922 347758 588222 347994
rect 588458 347758 588542 347994
rect 588778 347758 588810 347994
rect -4886 347576 588810 347758
rect -2966 344294 586890 344476
rect -2966 344058 -2934 344294
rect -2698 344058 -2614 344294
rect -2378 344058 18986 344294
rect 19222 344058 40328 344294
rect 40564 344058 176056 344294
rect 176292 344058 198986 344294
rect 199222 344058 234986 344294
rect 235222 344058 270986 344294
rect 271222 344058 306986 344294
rect 307222 344058 340328 344294
rect 340564 344058 476056 344294
rect 476292 344058 486986 344294
rect 487222 344058 522986 344294
rect 523222 344058 558986 344294
rect 559222 344058 586302 344294
rect 586538 344058 586622 344294
rect 586858 344058 586890 344294
rect -2966 343876 586890 344058
rect -8726 337394 592650 337576
rect -8726 337158 -7734 337394
rect -7498 337158 -7414 337394
rect -7178 337158 12086 337394
rect 12322 337158 48086 337394
rect 48322 337158 84086 337394
rect 84322 337158 120086 337394
rect 120322 337158 156086 337394
rect 156322 337158 192086 337394
rect 192322 337158 228086 337394
rect 228322 337158 264086 337394
rect 264322 337158 300086 337394
rect 300322 337158 336086 337394
rect 336322 337158 372086 337394
rect 372322 337158 408086 337394
rect 408322 337158 444086 337394
rect 444322 337158 480086 337394
rect 480322 337158 516086 337394
rect 516322 337158 552086 337394
rect 552322 337158 591102 337394
rect 591338 337158 591422 337394
rect 591658 337158 592650 337394
rect -8726 336976 592650 337158
rect -6806 333694 590730 333876
rect -6806 333458 -5814 333694
rect -5578 333458 -5494 333694
rect -5258 333458 8386 333694
rect 8622 333458 44386 333694
rect 44622 333458 80386 333694
rect 80622 333458 116386 333694
rect 116622 333458 152386 333694
rect 152622 333458 188386 333694
rect 188622 333458 224386 333694
rect 224622 333458 260386 333694
rect 260622 333458 296386 333694
rect 296622 333458 332386 333694
rect 332622 333458 368386 333694
rect 368622 333458 404386 333694
rect 404622 333458 440386 333694
rect 440622 333458 476386 333694
rect 476622 333458 512386 333694
rect 512622 333458 548386 333694
rect 548622 333458 589182 333694
rect 589418 333458 589502 333694
rect 589738 333458 590730 333694
rect -6806 333276 590730 333458
rect -4886 329994 588810 330176
rect -4886 329758 -3894 329994
rect -3658 329758 -3574 329994
rect -3338 329758 4686 329994
rect 4922 329758 40686 329994
rect 40922 329758 76686 329994
rect 76922 329758 112686 329994
rect 112922 329758 148686 329994
rect 148922 329758 184686 329994
rect 184922 329758 220686 329994
rect 220922 329758 256686 329994
rect 256922 329758 292686 329994
rect 292922 329758 328686 329994
rect 328922 329758 364686 329994
rect 364922 329758 400686 329994
rect 400922 329758 436686 329994
rect 436922 329758 472686 329994
rect 472922 329758 508686 329994
rect 508922 329758 544686 329994
rect 544922 329758 580686 329994
rect 580922 329758 587262 329994
rect 587498 329758 587582 329994
rect 587818 329758 588810 329994
rect -4886 329576 588810 329758
rect -2966 326294 586890 326476
rect -2966 326058 -1974 326294
rect -1738 326058 -1654 326294
rect -1418 326058 986 326294
rect 1222 326058 36986 326294
rect 37222 326058 72986 326294
rect 73222 326058 108986 326294
rect 109222 326058 144986 326294
rect 145222 326058 180986 326294
rect 181222 326058 216986 326294
rect 217222 326058 252986 326294
rect 253222 326058 288986 326294
rect 289222 326058 324986 326294
rect 325222 326058 360986 326294
rect 361222 326058 396986 326294
rect 397222 326058 432986 326294
rect 433222 326058 468986 326294
rect 469222 326058 504986 326294
rect 505222 326058 540986 326294
rect 541222 326058 576986 326294
rect 577222 326058 585342 326294
rect 585578 326058 585662 326294
rect 585898 326058 586890 326294
rect -2966 325876 586890 326058
rect -8726 319394 592650 319576
rect -8726 319158 -8694 319394
rect -8458 319158 -8374 319394
rect -8138 319158 30086 319394
rect 30322 319158 66086 319394
rect 66322 319158 102086 319394
rect 102322 319158 138086 319394
rect 138322 319158 174086 319394
rect 174322 319158 210086 319394
rect 210322 319158 246086 319394
rect 246322 319158 282086 319394
rect 282322 319158 318086 319394
rect 318322 319158 354086 319394
rect 354322 319158 390086 319394
rect 390322 319158 426086 319394
rect 426322 319158 462086 319394
rect 462322 319158 498086 319394
rect 498322 319158 534086 319394
rect 534322 319158 570086 319394
rect 570322 319158 592062 319394
rect 592298 319158 592382 319394
rect 592618 319158 592650 319394
rect -8726 318976 592650 319158
rect -6806 315694 590730 315876
rect -6806 315458 -6774 315694
rect -6538 315458 -6454 315694
rect -6218 315458 26386 315694
rect 26622 315458 62386 315694
rect 62622 315458 98386 315694
rect 98622 315458 134386 315694
rect 134622 315458 170386 315694
rect 170622 315458 206386 315694
rect 206622 315458 242386 315694
rect 242622 315458 278386 315694
rect 278622 315458 314386 315694
rect 314622 315458 350386 315694
rect 350622 315458 386386 315694
rect 386622 315458 422386 315694
rect 422622 315458 458386 315694
rect 458622 315458 494386 315694
rect 494622 315458 530386 315694
rect 530622 315458 566386 315694
rect 566622 315458 590142 315694
rect 590378 315458 590462 315694
rect 590698 315458 590730 315694
rect -6806 315276 590730 315458
rect -4886 311994 588810 312176
rect -4886 311758 -4854 311994
rect -4618 311758 -4534 311994
rect -4298 311758 22686 311994
rect 22922 311758 58686 311994
rect 58922 311758 94686 311994
rect 94922 311758 130686 311994
rect 130922 311758 166686 311994
rect 166922 311758 202686 311994
rect 202922 311758 238686 311994
rect 238922 311758 274686 311994
rect 274922 311758 310686 311994
rect 310922 311758 346686 311994
rect 346922 311758 382686 311994
rect 382922 311758 418686 311994
rect 418922 311758 454686 311994
rect 454922 311758 490686 311994
rect 490922 311758 526686 311994
rect 526922 311758 562686 311994
rect 562922 311758 588222 311994
rect 588458 311758 588542 311994
rect 588778 311758 588810 311994
rect -4886 311576 588810 311758
rect -2966 308294 586890 308476
rect -2966 308058 -2934 308294
rect -2698 308058 -2614 308294
rect -2378 308058 18986 308294
rect 19222 308058 54986 308294
rect 55222 308058 90986 308294
rect 91222 308058 126986 308294
rect 127222 308058 162986 308294
rect 163222 308058 198986 308294
rect 199222 308058 234986 308294
rect 235222 308058 270986 308294
rect 271222 308058 306986 308294
rect 307222 308058 342986 308294
rect 343222 308058 378986 308294
rect 379222 308058 414986 308294
rect 415222 308058 450986 308294
rect 451222 308058 486986 308294
rect 487222 308058 522986 308294
rect 523222 308058 558986 308294
rect 559222 308058 586302 308294
rect 586538 308058 586622 308294
rect 586858 308058 586890 308294
rect -2966 307876 586890 308058
rect -8726 301394 592650 301576
rect -8726 301158 -7734 301394
rect -7498 301158 -7414 301394
rect -7178 301158 12086 301394
rect 12322 301158 48086 301394
rect 48322 301158 84086 301394
rect 84322 301158 120086 301394
rect 120322 301158 156086 301394
rect 156322 301158 192086 301394
rect 192322 301158 228086 301394
rect 228322 301158 264086 301394
rect 264322 301158 300086 301394
rect 300322 301158 336086 301394
rect 336322 301158 372086 301394
rect 372322 301158 408086 301394
rect 408322 301158 444086 301394
rect 444322 301158 480086 301394
rect 480322 301158 516086 301394
rect 516322 301158 552086 301394
rect 552322 301158 591102 301394
rect 591338 301158 591422 301394
rect 591658 301158 592650 301394
rect -8726 300976 592650 301158
rect -6806 297694 590730 297876
rect -6806 297458 -5814 297694
rect -5578 297458 -5494 297694
rect -5258 297458 8386 297694
rect 8622 297458 44386 297694
rect 44622 297458 80386 297694
rect 80622 297458 116386 297694
rect 116622 297458 152386 297694
rect 152622 297458 188386 297694
rect 188622 297458 224386 297694
rect 224622 297458 260386 297694
rect 260622 297458 296386 297694
rect 296622 297458 332386 297694
rect 332622 297458 368386 297694
rect 368622 297458 404386 297694
rect 404622 297458 440386 297694
rect 440622 297458 476386 297694
rect 476622 297458 512386 297694
rect 512622 297458 548386 297694
rect 548622 297458 589182 297694
rect 589418 297458 589502 297694
rect 589738 297458 590730 297694
rect -6806 297276 590730 297458
rect -4886 293994 588810 294176
rect -4886 293758 -3894 293994
rect -3658 293758 -3574 293994
rect -3338 293758 4686 293994
rect 4922 293758 40686 293994
rect 40922 293758 76686 293994
rect 76922 293758 112686 293994
rect 112922 293758 148686 293994
rect 148922 293758 184686 293994
rect 184922 293758 220686 293994
rect 220922 293758 256686 293994
rect 256922 293758 292686 293994
rect 292922 293758 328686 293994
rect 328922 293758 364686 293994
rect 364922 293758 400686 293994
rect 400922 293758 436686 293994
rect 436922 293758 472686 293994
rect 472922 293758 508686 293994
rect 508922 293758 544686 293994
rect 544922 293758 580686 293994
rect 580922 293758 587262 293994
rect 587498 293758 587582 293994
rect 587818 293758 588810 293994
rect -4886 293576 588810 293758
rect -2966 290294 586890 290476
rect -2966 290058 -1974 290294
rect -1738 290058 -1654 290294
rect -1418 290058 986 290294
rect 1222 290058 36986 290294
rect 37222 290058 72986 290294
rect 73222 290058 108986 290294
rect 109222 290058 144986 290294
rect 145222 290058 180986 290294
rect 181222 290058 216986 290294
rect 217222 290058 252986 290294
rect 253222 290058 288986 290294
rect 289222 290058 324986 290294
rect 325222 290058 360986 290294
rect 361222 290058 396986 290294
rect 397222 290058 432986 290294
rect 433222 290058 468986 290294
rect 469222 290058 504986 290294
rect 505222 290058 540986 290294
rect 541222 290058 576986 290294
rect 577222 290058 585342 290294
rect 585578 290058 585662 290294
rect 585898 290058 586890 290294
rect -2966 289876 586890 290058
rect -8726 283394 592650 283576
rect -8726 283158 -8694 283394
rect -8458 283158 -8374 283394
rect -8138 283158 30086 283394
rect 30322 283158 66086 283394
rect 66322 283158 102086 283394
rect 102322 283158 138086 283394
rect 138322 283158 174086 283394
rect 174322 283158 210086 283394
rect 210322 283158 246086 283394
rect 246322 283158 282086 283394
rect 282322 283158 318086 283394
rect 318322 283158 354086 283394
rect 354322 283158 390086 283394
rect 390322 283158 426086 283394
rect 426322 283158 462086 283394
rect 462322 283158 498086 283394
rect 498322 283158 534086 283394
rect 534322 283158 570086 283394
rect 570322 283158 592062 283394
rect 592298 283158 592382 283394
rect 592618 283158 592650 283394
rect -8726 282976 592650 283158
rect -6806 279694 590730 279876
rect -6806 279458 -6774 279694
rect -6538 279458 -6454 279694
rect -6218 279458 26386 279694
rect 26622 279458 62386 279694
rect 62622 279458 98386 279694
rect 98622 279458 134386 279694
rect 134622 279458 170386 279694
rect 170622 279458 206386 279694
rect 206622 279458 242386 279694
rect 242622 279458 278386 279694
rect 278622 279458 314386 279694
rect 314622 279458 350386 279694
rect 350622 279458 386386 279694
rect 386622 279458 422386 279694
rect 422622 279458 458386 279694
rect 458622 279458 494386 279694
rect 494622 279458 530386 279694
rect 530622 279458 566386 279694
rect 566622 279458 590142 279694
rect 590378 279458 590462 279694
rect 590698 279458 590730 279694
rect -6806 279276 590730 279458
rect -4886 275994 588810 276176
rect -4886 275758 -4854 275994
rect -4618 275758 -4534 275994
rect -4298 275758 22686 275994
rect 22922 275758 58686 275994
rect 58922 275758 94686 275994
rect 94922 275758 130686 275994
rect 130922 275758 166686 275994
rect 166922 275758 202686 275994
rect 202922 275758 238686 275994
rect 238922 275758 274686 275994
rect 274922 275758 310686 275994
rect 310922 275758 346686 275994
rect 346922 275758 382686 275994
rect 382922 275758 418686 275994
rect 418922 275758 454686 275994
rect 454922 275758 490686 275994
rect 490922 275758 526686 275994
rect 526922 275758 562686 275994
rect 562922 275758 588222 275994
rect 588458 275758 588542 275994
rect 588778 275758 588810 275994
rect -4886 275576 588810 275758
rect -2966 272294 586890 272476
rect -2966 272058 -2934 272294
rect -2698 272058 -2614 272294
rect -2378 272058 18986 272294
rect 19222 272058 54986 272294
rect 55222 272058 90986 272294
rect 91222 272058 126986 272294
rect 127222 272058 162986 272294
rect 163222 272058 198986 272294
rect 199222 272058 234986 272294
rect 235222 272058 270986 272294
rect 271222 272058 306986 272294
rect 307222 272058 342986 272294
rect 343222 272058 378986 272294
rect 379222 272058 414986 272294
rect 415222 272058 450986 272294
rect 451222 272058 486986 272294
rect 487222 272058 522986 272294
rect 523222 272058 558986 272294
rect 559222 272058 586302 272294
rect 586538 272058 586622 272294
rect 586858 272058 586890 272294
rect -2966 271876 586890 272058
rect -8726 265394 592650 265576
rect -8726 265158 -7734 265394
rect -7498 265158 -7414 265394
rect -7178 265158 12086 265394
rect 12322 265158 48086 265394
rect 48322 265158 84086 265394
rect 84322 265158 120086 265394
rect 120322 265158 156086 265394
rect 156322 265158 192086 265394
rect 192322 265158 228086 265394
rect 228322 265158 264086 265394
rect 264322 265158 300086 265394
rect 300322 265158 336086 265394
rect 336322 265158 372086 265394
rect 372322 265158 408086 265394
rect 408322 265158 444086 265394
rect 444322 265158 480086 265394
rect 480322 265158 516086 265394
rect 516322 265158 552086 265394
rect 552322 265158 591102 265394
rect 591338 265158 591422 265394
rect 591658 265158 592650 265394
rect -8726 264976 592650 265158
rect -6806 261694 590730 261876
rect -6806 261458 -5814 261694
rect -5578 261458 -5494 261694
rect -5258 261458 8386 261694
rect 8622 261458 44386 261694
rect 44622 261458 80386 261694
rect 80622 261458 116386 261694
rect 116622 261458 152386 261694
rect 152622 261458 188386 261694
rect 188622 261458 224386 261694
rect 224622 261458 260386 261694
rect 260622 261458 296386 261694
rect 296622 261458 332386 261694
rect 332622 261458 368386 261694
rect 368622 261458 404386 261694
rect 404622 261458 440386 261694
rect 440622 261458 476386 261694
rect 476622 261458 512386 261694
rect 512622 261458 548386 261694
rect 548622 261458 589182 261694
rect 589418 261458 589502 261694
rect 589738 261458 590730 261694
rect -6806 261276 590730 261458
rect -4886 257994 588810 258176
rect -4886 257758 -3894 257994
rect -3658 257758 -3574 257994
rect -3338 257758 4686 257994
rect 4922 257758 40686 257994
rect 40922 257758 76686 257994
rect 76922 257758 112686 257994
rect 112922 257758 148686 257994
rect 148922 257758 184686 257994
rect 184922 257758 220686 257994
rect 220922 257758 256686 257994
rect 256922 257758 292686 257994
rect 292922 257758 328686 257994
rect 328922 257758 364686 257994
rect 364922 257758 400686 257994
rect 400922 257758 436686 257994
rect 436922 257758 472686 257994
rect 472922 257758 508686 257994
rect 508922 257758 544686 257994
rect 544922 257758 580686 257994
rect 580922 257758 587262 257994
rect 587498 257758 587582 257994
rect 587818 257758 588810 257994
rect -4886 257576 588810 257758
rect -2966 254294 586890 254476
rect -2966 254058 -1974 254294
rect -1738 254058 -1654 254294
rect -1418 254058 986 254294
rect 1222 254058 36986 254294
rect 37222 254058 72986 254294
rect 73222 254058 108986 254294
rect 109222 254058 144986 254294
rect 145222 254058 180986 254294
rect 181222 254058 216986 254294
rect 217222 254058 252986 254294
rect 253222 254058 288986 254294
rect 289222 254058 324986 254294
rect 325222 254058 360986 254294
rect 361222 254058 396986 254294
rect 397222 254058 432986 254294
rect 433222 254058 468986 254294
rect 469222 254058 504986 254294
rect 505222 254058 540986 254294
rect 541222 254058 576986 254294
rect 577222 254058 585342 254294
rect 585578 254058 585662 254294
rect 585898 254058 586890 254294
rect -2966 253876 586890 254058
rect -8726 247394 592650 247576
rect -8726 247158 -8694 247394
rect -8458 247158 -8374 247394
rect -8138 247158 30086 247394
rect 30322 247158 66086 247394
rect 66322 247158 102086 247394
rect 102322 247158 138086 247394
rect 138322 247158 174086 247394
rect 174322 247158 210086 247394
rect 210322 247158 246086 247394
rect 246322 247158 282086 247394
rect 282322 247158 318086 247394
rect 318322 247158 354086 247394
rect 354322 247158 390086 247394
rect 390322 247158 426086 247394
rect 426322 247158 462086 247394
rect 462322 247158 498086 247394
rect 498322 247158 534086 247394
rect 534322 247158 570086 247394
rect 570322 247158 592062 247394
rect 592298 247158 592382 247394
rect 592618 247158 592650 247394
rect -8726 246976 592650 247158
rect -6806 243694 590730 243876
rect -6806 243458 -6774 243694
rect -6538 243458 -6454 243694
rect -6218 243458 26386 243694
rect 26622 243458 242386 243694
rect 242622 243458 278386 243694
rect 278622 243458 314386 243694
rect 314622 243458 350386 243694
rect 350622 243458 386386 243694
rect 386622 243458 422386 243694
rect 422622 243458 458386 243694
rect 458622 243458 494386 243694
rect 494622 243458 530386 243694
rect 530622 243458 566386 243694
rect 566622 243458 590142 243694
rect 590378 243458 590462 243694
rect 590698 243458 590730 243694
rect -6806 243276 590730 243458
rect -4886 239994 588810 240176
rect -4886 239758 -4854 239994
rect -4618 239758 -4534 239994
rect -4298 239758 22686 239994
rect 22922 239758 274686 239994
rect 274922 239758 310686 239994
rect 310922 239758 346686 239994
rect 346922 239758 382686 239994
rect 382922 239758 418686 239994
rect 418922 239758 454686 239994
rect 454922 239758 490686 239994
rect 490922 239758 526686 239994
rect 526922 239758 562686 239994
rect 562922 239758 588222 239994
rect 588458 239758 588542 239994
rect 588778 239758 588810 239994
rect -4886 239576 588810 239758
rect -2966 236294 586890 236476
rect -2966 236058 -2934 236294
rect -2698 236058 -2614 236294
rect -2378 236058 18986 236294
rect 19222 236058 59610 236294
rect 59846 236058 90330 236294
rect 90566 236058 121050 236294
rect 121286 236058 151770 236294
rect 152006 236058 182490 236294
rect 182726 236058 213210 236294
rect 213446 236058 270986 236294
rect 271222 236058 306986 236294
rect 307222 236058 342986 236294
rect 343222 236058 378986 236294
rect 379222 236058 414986 236294
rect 415222 236058 450986 236294
rect 451222 236058 486986 236294
rect 487222 236058 522986 236294
rect 523222 236058 558986 236294
rect 559222 236058 586302 236294
rect 586538 236058 586622 236294
rect 586858 236058 586890 236294
rect -2966 235876 586890 236058
rect -8726 229394 592650 229576
rect -8726 229158 -7734 229394
rect -7498 229158 -7414 229394
rect -7178 229158 12086 229394
rect 12322 229158 264086 229394
rect 264322 229158 300086 229394
rect 300322 229158 336086 229394
rect 336322 229158 372086 229394
rect 372322 229158 408086 229394
rect 408322 229158 444086 229394
rect 444322 229158 480086 229394
rect 480322 229158 516086 229394
rect 516322 229158 552086 229394
rect 552322 229158 591102 229394
rect 591338 229158 591422 229394
rect 591658 229158 592650 229394
rect -8726 228976 592650 229158
rect -6806 225694 590730 225876
rect -6806 225458 -5814 225694
rect -5578 225458 -5494 225694
rect -5258 225458 8386 225694
rect 8622 225458 260386 225694
rect 260622 225458 296386 225694
rect 296622 225458 332386 225694
rect 332622 225458 368386 225694
rect 368622 225458 404386 225694
rect 404622 225458 440386 225694
rect 440622 225458 476386 225694
rect 476622 225458 512386 225694
rect 512622 225458 548386 225694
rect 548622 225458 589182 225694
rect 589418 225458 589502 225694
rect 589738 225458 590730 225694
rect -6806 225276 590730 225458
rect -4886 221994 588810 222176
rect -4886 221758 -3894 221994
rect -3658 221758 -3574 221994
rect -3338 221758 4686 221994
rect 4922 221758 256686 221994
rect 256922 221758 292686 221994
rect 292922 221758 328686 221994
rect 328922 221758 364686 221994
rect 364922 221758 400686 221994
rect 400922 221758 436686 221994
rect 436922 221758 472686 221994
rect 472922 221758 508686 221994
rect 508922 221758 544686 221994
rect 544922 221758 580686 221994
rect 580922 221758 587262 221994
rect 587498 221758 587582 221994
rect 587818 221758 588810 221994
rect -4886 221576 588810 221758
rect -2966 218294 586890 218476
rect -2966 218058 -1974 218294
rect -1738 218058 -1654 218294
rect -1418 218058 986 218294
rect 1222 218058 36986 218294
rect 37222 218058 44250 218294
rect 44486 218058 74970 218294
rect 75206 218058 105690 218294
rect 105926 218058 136410 218294
rect 136646 218058 167130 218294
rect 167366 218058 197850 218294
rect 198086 218058 228570 218294
rect 228806 218058 252986 218294
rect 253222 218058 288986 218294
rect 289222 218058 324986 218294
rect 325222 218058 360986 218294
rect 361222 218058 396986 218294
rect 397222 218058 432986 218294
rect 433222 218058 468986 218294
rect 469222 218058 504986 218294
rect 505222 218058 540986 218294
rect 541222 218058 576986 218294
rect 577222 218058 585342 218294
rect 585578 218058 585662 218294
rect 585898 218058 586890 218294
rect -2966 217876 586890 218058
rect -8726 211394 592650 211576
rect -8726 211158 -8694 211394
rect -8458 211158 -8374 211394
rect -8138 211158 30086 211394
rect 30322 211158 246086 211394
rect 246322 211158 282086 211394
rect 282322 211158 318086 211394
rect 318322 211158 354086 211394
rect 354322 211158 390086 211394
rect 390322 211158 426086 211394
rect 426322 211158 462086 211394
rect 462322 211158 498086 211394
rect 498322 211158 534086 211394
rect 534322 211158 570086 211394
rect 570322 211158 592062 211394
rect 592298 211158 592382 211394
rect 592618 211158 592650 211394
rect -8726 210976 592650 211158
rect -6806 207694 590730 207876
rect -6806 207458 -6774 207694
rect -6538 207458 -6454 207694
rect -6218 207458 26386 207694
rect 26622 207458 242386 207694
rect 242622 207458 278386 207694
rect 278622 207458 314386 207694
rect 314622 207458 350386 207694
rect 350622 207458 386386 207694
rect 386622 207458 422386 207694
rect 422622 207458 458386 207694
rect 458622 207458 494386 207694
rect 494622 207458 530386 207694
rect 530622 207458 566386 207694
rect 566622 207458 590142 207694
rect 590378 207458 590462 207694
rect 590698 207458 590730 207694
rect -6806 207276 590730 207458
rect -4886 203994 588810 204176
rect -4886 203758 -4854 203994
rect -4618 203758 -4534 203994
rect -4298 203758 22686 203994
rect 22922 203758 274686 203994
rect 274922 203758 310686 203994
rect 310922 203758 346686 203994
rect 346922 203758 382686 203994
rect 382922 203758 418686 203994
rect 418922 203758 454686 203994
rect 454922 203758 490686 203994
rect 490922 203758 526686 203994
rect 526922 203758 562686 203994
rect 562922 203758 588222 203994
rect 588458 203758 588542 203994
rect 588778 203758 588810 203994
rect -4886 203576 588810 203758
rect -2966 200294 586890 200476
rect -2966 200058 -2934 200294
rect -2698 200058 -2614 200294
rect -2378 200058 18986 200294
rect 19222 200058 59610 200294
rect 59846 200058 90330 200294
rect 90566 200058 121050 200294
rect 121286 200058 151770 200294
rect 152006 200058 182490 200294
rect 182726 200058 213210 200294
rect 213446 200058 270986 200294
rect 271222 200058 306986 200294
rect 307222 200058 342986 200294
rect 343222 200058 378986 200294
rect 379222 200058 414986 200294
rect 415222 200058 450986 200294
rect 451222 200058 486986 200294
rect 487222 200058 522986 200294
rect 523222 200058 558986 200294
rect 559222 200058 586302 200294
rect 586538 200058 586622 200294
rect 586858 200058 586890 200294
rect -2966 199876 586890 200058
rect -8726 193394 592650 193576
rect -8726 193158 -7734 193394
rect -7498 193158 -7414 193394
rect -7178 193158 12086 193394
rect 12322 193158 264086 193394
rect 264322 193158 300086 193394
rect 300322 193158 336086 193394
rect 336322 193158 372086 193394
rect 372322 193158 408086 193394
rect 408322 193158 444086 193394
rect 444322 193158 480086 193394
rect 480322 193158 516086 193394
rect 516322 193158 552086 193394
rect 552322 193158 591102 193394
rect 591338 193158 591422 193394
rect 591658 193158 592650 193394
rect -8726 192976 592650 193158
rect -6806 189694 590730 189876
rect -6806 189458 -5814 189694
rect -5578 189458 -5494 189694
rect -5258 189458 8386 189694
rect 8622 189458 260386 189694
rect 260622 189458 296386 189694
rect 296622 189458 332386 189694
rect 332622 189458 368386 189694
rect 368622 189458 404386 189694
rect 404622 189458 440386 189694
rect 440622 189458 476386 189694
rect 476622 189458 512386 189694
rect 512622 189458 548386 189694
rect 548622 189458 589182 189694
rect 589418 189458 589502 189694
rect 589738 189458 590730 189694
rect -6806 189276 590730 189458
rect -4886 185994 588810 186176
rect -4886 185758 -3894 185994
rect -3658 185758 -3574 185994
rect -3338 185758 4686 185994
rect 4922 185758 256686 185994
rect 256922 185758 292686 185994
rect 292922 185758 328686 185994
rect 328922 185758 364686 185994
rect 364922 185758 400686 185994
rect 400922 185758 436686 185994
rect 436922 185758 472686 185994
rect 472922 185758 508686 185994
rect 508922 185758 544686 185994
rect 544922 185758 580686 185994
rect 580922 185758 587262 185994
rect 587498 185758 587582 185994
rect 587818 185758 588810 185994
rect -4886 185576 588810 185758
rect -2966 182294 586890 182476
rect -2966 182058 -1974 182294
rect -1738 182058 -1654 182294
rect -1418 182058 986 182294
rect 1222 182058 36986 182294
rect 37222 182058 44250 182294
rect 44486 182058 74970 182294
rect 75206 182058 105690 182294
rect 105926 182058 136410 182294
rect 136646 182058 167130 182294
rect 167366 182058 197850 182294
rect 198086 182058 228570 182294
rect 228806 182058 252986 182294
rect 253222 182058 288986 182294
rect 289222 182058 324986 182294
rect 325222 182058 360986 182294
rect 361222 182058 396986 182294
rect 397222 182058 432986 182294
rect 433222 182058 468986 182294
rect 469222 182058 504986 182294
rect 505222 182058 540986 182294
rect 541222 182058 576986 182294
rect 577222 182058 585342 182294
rect 585578 182058 585662 182294
rect 585898 182058 586890 182294
rect -2966 181876 586890 182058
rect -8726 175394 592650 175576
rect -8726 175158 -8694 175394
rect -8458 175158 -8374 175394
rect -8138 175158 30086 175394
rect 30322 175158 246086 175394
rect 246322 175158 282086 175394
rect 282322 175158 318086 175394
rect 318322 175158 354086 175394
rect 354322 175158 390086 175394
rect 390322 175158 426086 175394
rect 426322 175158 462086 175394
rect 462322 175158 498086 175394
rect 498322 175158 534086 175394
rect 534322 175158 570086 175394
rect 570322 175158 592062 175394
rect 592298 175158 592382 175394
rect 592618 175158 592650 175394
rect -8726 174976 592650 175158
rect -6806 171694 590730 171876
rect -6806 171458 -6774 171694
rect -6538 171458 -6454 171694
rect -6218 171458 26386 171694
rect 26622 171458 242386 171694
rect 242622 171458 278386 171694
rect 278622 171458 314386 171694
rect 314622 171458 350386 171694
rect 350622 171458 386386 171694
rect 386622 171458 422386 171694
rect 422622 171458 458386 171694
rect 458622 171458 494386 171694
rect 494622 171458 530386 171694
rect 530622 171458 566386 171694
rect 566622 171458 590142 171694
rect 590378 171458 590462 171694
rect 590698 171458 590730 171694
rect -6806 171276 590730 171458
rect -4886 167994 588810 168176
rect -4886 167758 -4854 167994
rect -4618 167758 -4534 167994
rect -4298 167758 22686 167994
rect 22922 167758 274686 167994
rect 274922 167758 310686 167994
rect 310922 167758 346686 167994
rect 346922 167758 382686 167994
rect 382922 167758 418686 167994
rect 418922 167758 454686 167994
rect 454922 167758 490686 167994
rect 490922 167758 526686 167994
rect 526922 167758 562686 167994
rect 562922 167758 588222 167994
rect 588458 167758 588542 167994
rect 588778 167758 588810 167994
rect -4886 167576 588810 167758
rect -2966 164294 586890 164476
rect -2966 164058 -2934 164294
rect -2698 164058 -2614 164294
rect -2378 164058 18986 164294
rect 19222 164058 59610 164294
rect 59846 164058 90330 164294
rect 90566 164058 121050 164294
rect 121286 164058 151770 164294
rect 152006 164058 182490 164294
rect 182726 164058 213210 164294
rect 213446 164058 270986 164294
rect 271222 164058 306986 164294
rect 307222 164058 342986 164294
rect 343222 164058 378986 164294
rect 379222 164058 414986 164294
rect 415222 164058 450986 164294
rect 451222 164058 486986 164294
rect 487222 164058 522986 164294
rect 523222 164058 558986 164294
rect 559222 164058 586302 164294
rect 586538 164058 586622 164294
rect 586858 164058 586890 164294
rect -2966 163876 586890 164058
rect -8726 157394 592650 157576
rect -8726 157158 -7734 157394
rect -7498 157158 -7414 157394
rect -7178 157158 12086 157394
rect 12322 157158 264086 157394
rect 264322 157158 300086 157394
rect 300322 157158 336086 157394
rect 336322 157158 372086 157394
rect 372322 157158 408086 157394
rect 408322 157158 444086 157394
rect 444322 157158 480086 157394
rect 480322 157158 516086 157394
rect 516322 157158 552086 157394
rect 552322 157158 591102 157394
rect 591338 157158 591422 157394
rect 591658 157158 592650 157394
rect -8726 156976 592650 157158
rect -6806 153694 590730 153876
rect -6806 153458 -5814 153694
rect -5578 153458 -5494 153694
rect -5258 153458 8386 153694
rect 8622 153458 260386 153694
rect 260622 153458 296386 153694
rect 296622 153458 332386 153694
rect 332622 153458 368386 153694
rect 368622 153458 404386 153694
rect 404622 153458 440386 153694
rect 440622 153458 476386 153694
rect 476622 153458 512386 153694
rect 512622 153458 548386 153694
rect 548622 153458 589182 153694
rect 589418 153458 589502 153694
rect 589738 153458 590730 153694
rect -6806 153276 590730 153458
rect -4886 149994 588810 150176
rect -4886 149758 -3894 149994
rect -3658 149758 -3574 149994
rect -3338 149758 4686 149994
rect 4922 149758 256686 149994
rect 256922 149758 292686 149994
rect 292922 149758 328686 149994
rect 328922 149758 364686 149994
rect 364922 149758 400686 149994
rect 400922 149758 436686 149994
rect 436922 149758 472686 149994
rect 472922 149758 508686 149994
rect 508922 149758 544686 149994
rect 544922 149758 580686 149994
rect 580922 149758 587262 149994
rect 587498 149758 587582 149994
rect 587818 149758 588810 149994
rect -4886 149576 588810 149758
rect -2966 146294 586890 146476
rect -2966 146058 -1974 146294
rect -1738 146058 -1654 146294
rect -1418 146058 986 146294
rect 1222 146058 36986 146294
rect 37222 146058 44250 146294
rect 44486 146058 74970 146294
rect 75206 146058 105690 146294
rect 105926 146058 136410 146294
rect 136646 146058 167130 146294
rect 167366 146058 197850 146294
rect 198086 146058 228570 146294
rect 228806 146058 252986 146294
rect 253222 146058 288986 146294
rect 289222 146058 324986 146294
rect 325222 146058 360986 146294
rect 361222 146058 396986 146294
rect 397222 146058 432986 146294
rect 433222 146058 468986 146294
rect 469222 146058 504986 146294
rect 505222 146058 540986 146294
rect 541222 146058 576986 146294
rect 577222 146058 585342 146294
rect 585578 146058 585662 146294
rect 585898 146058 586890 146294
rect -2966 145876 586890 146058
rect -8726 139394 592650 139576
rect -8726 139158 -8694 139394
rect -8458 139158 -8374 139394
rect -8138 139158 30086 139394
rect 30322 139158 246086 139394
rect 246322 139158 282086 139394
rect 282322 139158 318086 139394
rect 318322 139158 354086 139394
rect 354322 139158 390086 139394
rect 390322 139158 426086 139394
rect 426322 139158 462086 139394
rect 462322 139158 498086 139394
rect 498322 139158 534086 139394
rect 534322 139158 570086 139394
rect 570322 139158 592062 139394
rect 592298 139158 592382 139394
rect 592618 139158 592650 139394
rect -8726 138976 592650 139158
rect -6806 135694 590730 135876
rect -6806 135458 -6774 135694
rect -6538 135458 -6454 135694
rect -6218 135458 26386 135694
rect 26622 135458 242386 135694
rect 242622 135458 278386 135694
rect 278622 135458 314386 135694
rect 314622 135458 350386 135694
rect 350622 135458 386386 135694
rect 386622 135458 422386 135694
rect 422622 135458 458386 135694
rect 458622 135458 494386 135694
rect 494622 135458 530386 135694
rect 530622 135458 566386 135694
rect 566622 135458 590142 135694
rect 590378 135458 590462 135694
rect 590698 135458 590730 135694
rect -6806 135276 590730 135458
rect -4886 131994 588810 132176
rect -4886 131758 -4854 131994
rect -4618 131758 -4534 131994
rect -4298 131758 22686 131994
rect 22922 131758 274686 131994
rect 274922 131758 310686 131994
rect 310922 131758 346686 131994
rect 346922 131758 382686 131994
rect 382922 131758 418686 131994
rect 418922 131758 454686 131994
rect 454922 131758 490686 131994
rect 490922 131758 526686 131994
rect 526922 131758 562686 131994
rect 562922 131758 588222 131994
rect 588458 131758 588542 131994
rect 588778 131758 588810 131994
rect -4886 131576 588810 131758
rect -2966 128294 586890 128476
rect -2966 128058 -2934 128294
rect -2698 128058 -2614 128294
rect -2378 128058 18986 128294
rect 19222 128058 59610 128294
rect 59846 128058 90330 128294
rect 90566 128058 121050 128294
rect 121286 128058 151770 128294
rect 152006 128058 182490 128294
rect 182726 128058 213210 128294
rect 213446 128058 270986 128294
rect 271222 128058 306986 128294
rect 307222 128058 342986 128294
rect 343222 128058 378986 128294
rect 379222 128058 414986 128294
rect 415222 128058 450986 128294
rect 451222 128058 486986 128294
rect 487222 128058 522986 128294
rect 523222 128058 558986 128294
rect 559222 128058 586302 128294
rect 586538 128058 586622 128294
rect 586858 128058 586890 128294
rect -2966 127876 586890 128058
rect -8726 121394 592650 121576
rect -8726 121158 -7734 121394
rect -7498 121158 -7414 121394
rect -7178 121158 12086 121394
rect 12322 121158 264086 121394
rect 264322 121158 300086 121394
rect 300322 121158 336086 121394
rect 336322 121158 372086 121394
rect 372322 121158 408086 121394
rect 408322 121158 444086 121394
rect 444322 121158 480086 121394
rect 480322 121158 516086 121394
rect 516322 121158 552086 121394
rect 552322 121158 591102 121394
rect 591338 121158 591422 121394
rect 591658 121158 592650 121394
rect -8726 120976 592650 121158
rect -6806 117694 590730 117876
rect -6806 117458 -5814 117694
rect -5578 117458 -5494 117694
rect -5258 117458 8386 117694
rect 8622 117458 260386 117694
rect 260622 117458 296386 117694
rect 296622 117458 332386 117694
rect 332622 117458 368386 117694
rect 368622 117458 404386 117694
rect 404622 117458 440386 117694
rect 440622 117458 476386 117694
rect 476622 117458 512386 117694
rect 512622 117458 548386 117694
rect 548622 117458 589182 117694
rect 589418 117458 589502 117694
rect 589738 117458 590730 117694
rect -6806 117276 590730 117458
rect -4886 113994 588810 114176
rect -4886 113758 -3894 113994
rect -3658 113758 -3574 113994
rect -3338 113758 4686 113994
rect 4922 113758 256686 113994
rect 256922 113758 292686 113994
rect 292922 113758 328686 113994
rect 328922 113758 364686 113994
rect 364922 113758 400686 113994
rect 400922 113758 436686 113994
rect 436922 113758 472686 113994
rect 472922 113758 508686 113994
rect 508922 113758 544686 113994
rect 544922 113758 580686 113994
rect 580922 113758 587262 113994
rect 587498 113758 587582 113994
rect 587818 113758 588810 113994
rect -4886 113576 588810 113758
rect -2966 110294 586890 110476
rect -2966 110058 -1974 110294
rect -1738 110058 -1654 110294
rect -1418 110058 986 110294
rect 1222 110058 36986 110294
rect 37222 110058 44250 110294
rect 44486 110058 74970 110294
rect 75206 110058 105690 110294
rect 105926 110058 136410 110294
rect 136646 110058 167130 110294
rect 167366 110058 197850 110294
rect 198086 110058 228570 110294
rect 228806 110058 252986 110294
rect 253222 110058 288986 110294
rect 289222 110058 324986 110294
rect 325222 110058 360986 110294
rect 361222 110058 396986 110294
rect 397222 110058 432986 110294
rect 433222 110058 468986 110294
rect 469222 110058 504986 110294
rect 505222 110058 540986 110294
rect 541222 110058 576986 110294
rect 577222 110058 585342 110294
rect 585578 110058 585662 110294
rect 585898 110058 586890 110294
rect -2966 109876 586890 110058
rect -8726 103394 592650 103576
rect -8726 103158 -8694 103394
rect -8458 103158 -8374 103394
rect -8138 103158 30086 103394
rect 30322 103158 246086 103394
rect 246322 103158 282086 103394
rect 282322 103158 318086 103394
rect 318322 103158 354086 103394
rect 354322 103158 390086 103394
rect 390322 103158 426086 103394
rect 426322 103158 462086 103394
rect 462322 103158 498086 103394
rect 498322 103158 534086 103394
rect 534322 103158 570086 103394
rect 570322 103158 592062 103394
rect 592298 103158 592382 103394
rect 592618 103158 592650 103394
rect -8726 102976 592650 103158
rect -6806 99694 590730 99876
rect -6806 99458 -6774 99694
rect -6538 99458 -6454 99694
rect -6218 99458 26386 99694
rect 26622 99458 242386 99694
rect 242622 99458 278386 99694
rect 278622 99458 314386 99694
rect 314622 99458 350386 99694
rect 350622 99458 386386 99694
rect 386622 99458 422386 99694
rect 422622 99458 458386 99694
rect 458622 99458 494386 99694
rect 494622 99458 530386 99694
rect 530622 99458 566386 99694
rect 566622 99458 590142 99694
rect 590378 99458 590462 99694
rect 590698 99458 590730 99694
rect -6806 99276 590730 99458
rect -4886 95994 588810 96176
rect -4886 95758 -4854 95994
rect -4618 95758 -4534 95994
rect -4298 95758 22686 95994
rect 22922 95758 274686 95994
rect 274922 95758 310686 95994
rect 310922 95758 346686 95994
rect 346922 95758 382686 95994
rect 382922 95758 418686 95994
rect 418922 95758 454686 95994
rect 454922 95758 490686 95994
rect 490922 95758 526686 95994
rect 526922 95758 562686 95994
rect 562922 95758 588222 95994
rect 588458 95758 588542 95994
rect 588778 95758 588810 95994
rect -4886 95576 588810 95758
rect -2966 92294 586890 92476
rect -2966 92058 -2934 92294
rect -2698 92058 -2614 92294
rect -2378 92058 18986 92294
rect 19222 92058 59610 92294
rect 59846 92058 90330 92294
rect 90566 92058 121050 92294
rect 121286 92058 151770 92294
rect 152006 92058 182490 92294
rect 182726 92058 213210 92294
rect 213446 92058 270986 92294
rect 271222 92058 306986 92294
rect 307222 92058 342986 92294
rect 343222 92058 378986 92294
rect 379222 92058 414986 92294
rect 415222 92058 450986 92294
rect 451222 92058 486986 92294
rect 487222 92058 522986 92294
rect 523222 92058 558986 92294
rect 559222 92058 586302 92294
rect 586538 92058 586622 92294
rect 586858 92058 586890 92294
rect -2966 91876 586890 92058
rect -8726 85394 592650 85576
rect -8726 85158 -7734 85394
rect -7498 85158 -7414 85394
rect -7178 85158 12086 85394
rect 12322 85158 264086 85394
rect 264322 85158 300086 85394
rect 300322 85158 336086 85394
rect 336322 85158 372086 85394
rect 372322 85158 408086 85394
rect 408322 85158 444086 85394
rect 444322 85158 480086 85394
rect 480322 85158 516086 85394
rect 516322 85158 552086 85394
rect 552322 85158 591102 85394
rect 591338 85158 591422 85394
rect 591658 85158 592650 85394
rect -8726 84976 592650 85158
rect -6806 81694 590730 81876
rect -6806 81458 -5814 81694
rect -5578 81458 -5494 81694
rect -5258 81458 8386 81694
rect 8622 81458 260386 81694
rect 260622 81458 296386 81694
rect 296622 81458 332386 81694
rect 332622 81458 368386 81694
rect 368622 81458 404386 81694
rect 404622 81458 440386 81694
rect 440622 81458 476386 81694
rect 476622 81458 512386 81694
rect 512622 81458 548386 81694
rect 548622 81458 589182 81694
rect 589418 81458 589502 81694
rect 589738 81458 590730 81694
rect -6806 81276 590730 81458
rect -4886 77994 588810 78176
rect -4886 77758 -3894 77994
rect -3658 77758 -3574 77994
rect -3338 77758 4686 77994
rect 4922 77758 256686 77994
rect 256922 77758 292686 77994
rect 292922 77758 328686 77994
rect 328922 77758 364686 77994
rect 364922 77758 400686 77994
rect 400922 77758 436686 77994
rect 436922 77758 472686 77994
rect 472922 77758 508686 77994
rect 508922 77758 544686 77994
rect 544922 77758 580686 77994
rect 580922 77758 587262 77994
rect 587498 77758 587582 77994
rect 587818 77758 588810 77994
rect -4886 77576 588810 77758
rect -2966 74294 586890 74476
rect -2966 74058 -1974 74294
rect -1738 74058 -1654 74294
rect -1418 74058 986 74294
rect 1222 74058 36986 74294
rect 37222 74058 44250 74294
rect 44486 74058 74970 74294
rect 75206 74058 105690 74294
rect 105926 74058 136410 74294
rect 136646 74058 167130 74294
rect 167366 74058 197850 74294
rect 198086 74058 228570 74294
rect 228806 74058 252986 74294
rect 253222 74058 288986 74294
rect 289222 74058 324986 74294
rect 325222 74058 360986 74294
rect 361222 74058 396986 74294
rect 397222 74058 432986 74294
rect 433222 74058 468986 74294
rect 469222 74058 504986 74294
rect 505222 74058 540986 74294
rect 541222 74058 576986 74294
rect 577222 74058 585342 74294
rect 585578 74058 585662 74294
rect 585898 74058 586890 74294
rect -2966 73876 586890 74058
rect -8726 67394 592650 67576
rect -8726 67158 -8694 67394
rect -8458 67158 -8374 67394
rect -8138 67158 30086 67394
rect 30322 67158 246086 67394
rect 246322 67158 282086 67394
rect 282322 67158 318086 67394
rect 318322 67158 354086 67394
rect 354322 67158 390086 67394
rect 390322 67158 426086 67394
rect 426322 67158 462086 67394
rect 462322 67158 498086 67394
rect 498322 67158 534086 67394
rect 534322 67158 570086 67394
rect 570322 67158 592062 67394
rect 592298 67158 592382 67394
rect 592618 67158 592650 67394
rect -8726 66976 592650 67158
rect -6806 63694 590730 63876
rect -6806 63458 -6774 63694
rect -6538 63458 -6454 63694
rect -6218 63458 26386 63694
rect 26622 63458 242386 63694
rect 242622 63458 278386 63694
rect 278622 63458 314386 63694
rect 314622 63458 350386 63694
rect 350622 63458 386386 63694
rect 386622 63458 422386 63694
rect 422622 63458 458386 63694
rect 458622 63458 494386 63694
rect 494622 63458 530386 63694
rect 530622 63458 566386 63694
rect 566622 63458 590142 63694
rect 590378 63458 590462 63694
rect 590698 63458 590730 63694
rect -6806 63276 590730 63458
rect -4886 59994 588810 60176
rect -4886 59758 -4854 59994
rect -4618 59758 -4534 59994
rect -4298 59758 22686 59994
rect 22922 59758 274686 59994
rect 274922 59758 310686 59994
rect 310922 59758 346686 59994
rect 346922 59758 382686 59994
rect 382922 59758 418686 59994
rect 418922 59758 454686 59994
rect 454922 59758 490686 59994
rect 490922 59758 526686 59994
rect 526922 59758 562686 59994
rect 562922 59758 588222 59994
rect 588458 59758 588542 59994
rect 588778 59758 588810 59994
rect -4886 59576 588810 59758
rect -2966 56294 586890 56476
rect -2966 56058 -2934 56294
rect -2698 56058 -2614 56294
rect -2378 56058 18986 56294
rect 19222 56058 59610 56294
rect 59846 56058 90330 56294
rect 90566 56058 121050 56294
rect 121286 56058 151770 56294
rect 152006 56058 182490 56294
rect 182726 56058 213210 56294
rect 213446 56058 270986 56294
rect 271222 56058 306986 56294
rect 307222 56058 342986 56294
rect 343222 56058 378986 56294
rect 379222 56058 414986 56294
rect 415222 56058 450986 56294
rect 451222 56058 486986 56294
rect 487222 56058 522986 56294
rect 523222 56058 558986 56294
rect 559222 56058 586302 56294
rect 586538 56058 586622 56294
rect 586858 56058 586890 56294
rect -2966 55876 586890 56058
rect -8726 49394 592650 49576
rect -8726 49158 -7734 49394
rect -7498 49158 -7414 49394
rect -7178 49158 12086 49394
rect 12322 49158 264086 49394
rect 264322 49158 300086 49394
rect 300322 49158 336086 49394
rect 336322 49158 372086 49394
rect 372322 49158 408086 49394
rect 408322 49158 444086 49394
rect 444322 49158 480086 49394
rect 480322 49158 516086 49394
rect 516322 49158 552086 49394
rect 552322 49158 591102 49394
rect 591338 49158 591422 49394
rect 591658 49158 592650 49394
rect -8726 48976 592650 49158
rect -6806 45694 590730 45876
rect -6806 45458 -5814 45694
rect -5578 45458 -5494 45694
rect -5258 45458 8386 45694
rect 8622 45458 260386 45694
rect 260622 45458 296386 45694
rect 296622 45458 332386 45694
rect 332622 45458 368386 45694
rect 368622 45458 404386 45694
rect 404622 45458 440386 45694
rect 440622 45458 476386 45694
rect 476622 45458 512386 45694
rect 512622 45458 548386 45694
rect 548622 45458 589182 45694
rect 589418 45458 589502 45694
rect 589738 45458 590730 45694
rect -6806 45276 590730 45458
rect -4886 41994 588810 42176
rect -4886 41758 -3894 41994
rect -3658 41758 -3574 41994
rect -3338 41758 4686 41994
rect 4922 41758 256686 41994
rect 256922 41758 292686 41994
rect 292922 41758 328686 41994
rect 328922 41758 364686 41994
rect 364922 41758 400686 41994
rect 400922 41758 436686 41994
rect 436922 41758 472686 41994
rect 472922 41758 508686 41994
rect 508922 41758 544686 41994
rect 544922 41758 580686 41994
rect 580922 41758 587262 41994
rect 587498 41758 587582 41994
rect 587818 41758 588810 41994
rect -4886 41576 588810 41758
rect -2966 38294 586890 38476
rect -2966 38058 -1974 38294
rect -1738 38058 -1654 38294
rect -1418 38058 986 38294
rect 1222 38058 36986 38294
rect 37222 38058 252986 38294
rect 253222 38058 288986 38294
rect 289222 38058 324986 38294
rect 325222 38058 360986 38294
rect 361222 38058 396986 38294
rect 397222 38058 432986 38294
rect 433222 38058 468986 38294
rect 469222 38058 504986 38294
rect 505222 38058 540986 38294
rect 541222 38058 576986 38294
rect 577222 38058 585342 38294
rect 585578 38058 585662 38294
rect 585898 38058 586890 38294
rect -2966 37876 586890 38058
rect -8726 31394 592650 31576
rect -8726 31158 -8694 31394
rect -8458 31158 -8374 31394
rect -8138 31158 30086 31394
rect 30322 31158 66086 31394
rect 66322 31158 102086 31394
rect 102322 31158 138086 31394
rect 138322 31158 174086 31394
rect 174322 31158 210086 31394
rect 210322 31158 246086 31394
rect 246322 31158 282086 31394
rect 282322 31158 318086 31394
rect 318322 31158 354086 31394
rect 354322 31158 390086 31394
rect 390322 31158 426086 31394
rect 426322 31158 462086 31394
rect 462322 31158 498086 31394
rect 498322 31158 534086 31394
rect 534322 31158 570086 31394
rect 570322 31158 592062 31394
rect 592298 31158 592382 31394
rect 592618 31158 592650 31394
rect -8726 30976 592650 31158
rect -6806 27694 590730 27876
rect -6806 27458 -6774 27694
rect -6538 27458 -6454 27694
rect -6218 27458 26386 27694
rect 26622 27458 62386 27694
rect 62622 27458 98386 27694
rect 98622 27458 134386 27694
rect 134622 27458 170386 27694
rect 170622 27458 206386 27694
rect 206622 27458 242386 27694
rect 242622 27458 278386 27694
rect 278622 27458 314386 27694
rect 314622 27458 350386 27694
rect 350622 27458 386386 27694
rect 386622 27458 422386 27694
rect 422622 27458 458386 27694
rect 458622 27458 494386 27694
rect 494622 27458 530386 27694
rect 530622 27458 566386 27694
rect 566622 27458 590142 27694
rect 590378 27458 590462 27694
rect 590698 27458 590730 27694
rect -6806 27276 590730 27458
rect -4886 23994 588810 24176
rect -4886 23758 -4854 23994
rect -4618 23758 -4534 23994
rect -4298 23758 22686 23994
rect 22922 23758 58686 23994
rect 58922 23758 94686 23994
rect 94922 23758 130686 23994
rect 130922 23758 166686 23994
rect 166922 23758 202686 23994
rect 202922 23758 238686 23994
rect 238922 23758 274686 23994
rect 274922 23758 310686 23994
rect 310922 23758 346686 23994
rect 346922 23758 382686 23994
rect 382922 23758 418686 23994
rect 418922 23758 454686 23994
rect 454922 23758 490686 23994
rect 490922 23758 526686 23994
rect 526922 23758 562686 23994
rect 562922 23758 588222 23994
rect 588458 23758 588542 23994
rect 588778 23758 588810 23994
rect -4886 23576 588810 23758
rect -2966 20294 586890 20476
rect -2966 20058 -2934 20294
rect -2698 20058 -2614 20294
rect -2378 20058 18986 20294
rect 19222 20058 54986 20294
rect 55222 20058 90986 20294
rect 91222 20058 126986 20294
rect 127222 20058 162986 20294
rect 163222 20058 198986 20294
rect 199222 20058 234986 20294
rect 235222 20058 270986 20294
rect 271222 20058 306986 20294
rect 307222 20058 342986 20294
rect 343222 20058 378986 20294
rect 379222 20058 414986 20294
rect 415222 20058 450986 20294
rect 451222 20058 486986 20294
rect 487222 20058 522986 20294
rect 523222 20058 558986 20294
rect 559222 20058 586302 20294
rect 586538 20058 586622 20294
rect 586858 20058 586890 20294
rect -2966 19876 586890 20058
rect -8726 13394 592650 13576
rect -8726 13158 -7734 13394
rect -7498 13158 -7414 13394
rect -7178 13158 12086 13394
rect 12322 13158 48086 13394
rect 48322 13158 84086 13394
rect 84322 13158 120086 13394
rect 120322 13158 156086 13394
rect 156322 13158 192086 13394
rect 192322 13158 228086 13394
rect 228322 13158 264086 13394
rect 264322 13158 300086 13394
rect 300322 13158 336086 13394
rect 336322 13158 372086 13394
rect 372322 13158 408086 13394
rect 408322 13158 444086 13394
rect 444322 13158 480086 13394
rect 480322 13158 516086 13394
rect 516322 13158 552086 13394
rect 552322 13158 591102 13394
rect 591338 13158 591422 13394
rect 591658 13158 592650 13394
rect -8726 12976 592650 13158
rect -6806 9694 590730 9876
rect -6806 9458 -5814 9694
rect -5578 9458 -5494 9694
rect -5258 9458 8386 9694
rect 8622 9458 44386 9694
rect 44622 9458 80386 9694
rect 80622 9458 116386 9694
rect 116622 9458 152386 9694
rect 152622 9458 188386 9694
rect 188622 9458 224386 9694
rect 224622 9458 260386 9694
rect 260622 9458 296386 9694
rect 296622 9458 332386 9694
rect 332622 9458 368386 9694
rect 368622 9458 404386 9694
rect 404622 9458 440386 9694
rect 440622 9458 476386 9694
rect 476622 9458 512386 9694
rect 512622 9458 548386 9694
rect 548622 9458 589182 9694
rect 589418 9458 589502 9694
rect 589738 9458 590730 9694
rect -6806 9276 590730 9458
rect -4886 5994 588810 6176
rect -4886 5758 -3894 5994
rect -3658 5758 -3574 5994
rect -3338 5758 4686 5994
rect 4922 5758 40686 5994
rect 40922 5758 76686 5994
rect 76922 5758 112686 5994
rect 112922 5758 148686 5994
rect 148922 5758 184686 5994
rect 184922 5758 220686 5994
rect 220922 5758 256686 5994
rect 256922 5758 292686 5994
rect 292922 5758 328686 5994
rect 328922 5758 364686 5994
rect 364922 5758 400686 5994
rect 400922 5758 436686 5994
rect 436922 5758 472686 5994
rect 472922 5758 508686 5994
rect 508922 5758 544686 5994
rect 544922 5758 580686 5994
rect 580922 5758 587262 5994
rect 587498 5758 587582 5994
rect 587818 5758 588810 5994
rect -4886 5576 588810 5758
rect -2966 2294 586890 2476
rect -2966 2058 -1974 2294
rect -1738 2058 -1654 2294
rect -1418 2058 986 2294
rect 1222 2058 36986 2294
rect 37222 2058 72986 2294
rect 73222 2058 108986 2294
rect 109222 2058 144986 2294
rect 145222 2058 180986 2294
rect 181222 2058 216986 2294
rect 217222 2058 252986 2294
rect 253222 2058 288986 2294
rect 289222 2058 324986 2294
rect 325222 2058 360986 2294
rect 361222 2058 396986 2294
rect 397222 2058 432986 2294
rect 433222 2058 468986 2294
rect 469222 2058 504986 2294
rect 505222 2058 540986 2294
rect 541222 2058 576986 2294
rect 577222 2058 585342 2294
rect 585578 2058 585662 2294
rect 585898 2058 586890 2294
rect -2966 1876 586890 2058
rect -2006 -346 585930 -314
rect -2006 -582 -1974 -346
rect -1738 -582 -1654 -346
rect -1418 -582 986 -346
rect 1222 -582 36986 -346
rect 37222 -582 72986 -346
rect 73222 -582 108986 -346
rect 109222 -582 144986 -346
rect 145222 -582 180986 -346
rect 181222 -582 216986 -346
rect 217222 -582 252986 -346
rect 253222 -582 288986 -346
rect 289222 -582 324986 -346
rect 325222 -582 360986 -346
rect 361222 -582 396986 -346
rect 397222 -582 432986 -346
rect 433222 -582 468986 -346
rect 469222 -582 504986 -346
rect 505222 -582 540986 -346
rect 541222 -582 576986 -346
rect 577222 -582 585342 -346
rect 585578 -582 585662 -346
rect 585898 -582 585930 -346
rect -2006 -666 585930 -582
rect -2006 -902 -1974 -666
rect -1738 -902 -1654 -666
rect -1418 -902 986 -666
rect 1222 -902 36986 -666
rect 37222 -902 72986 -666
rect 73222 -902 108986 -666
rect 109222 -902 144986 -666
rect 145222 -902 180986 -666
rect 181222 -902 216986 -666
rect 217222 -902 252986 -666
rect 253222 -902 288986 -666
rect 289222 -902 324986 -666
rect 325222 -902 360986 -666
rect 361222 -902 396986 -666
rect 397222 -902 432986 -666
rect 433222 -902 468986 -666
rect 469222 -902 504986 -666
rect 505222 -902 540986 -666
rect 541222 -902 576986 -666
rect 577222 -902 585342 -666
rect 585578 -902 585662 -666
rect 585898 -902 585930 -666
rect -2006 -934 585930 -902
rect -2966 -1306 586890 -1274
rect -2966 -1542 -2934 -1306
rect -2698 -1542 -2614 -1306
rect -2378 -1542 18986 -1306
rect 19222 -1542 54986 -1306
rect 55222 -1542 90986 -1306
rect 91222 -1542 126986 -1306
rect 127222 -1542 162986 -1306
rect 163222 -1542 198986 -1306
rect 199222 -1542 234986 -1306
rect 235222 -1542 270986 -1306
rect 271222 -1542 306986 -1306
rect 307222 -1542 342986 -1306
rect 343222 -1542 378986 -1306
rect 379222 -1542 414986 -1306
rect 415222 -1542 450986 -1306
rect 451222 -1542 486986 -1306
rect 487222 -1542 522986 -1306
rect 523222 -1542 558986 -1306
rect 559222 -1542 586302 -1306
rect 586538 -1542 586622 -1306
rect 586858 -1542 586890 -1306
rect -2966 -1626 586890 -1542
rect -2966 -1862 -2934 -1626
rect -2698 -1862 -2614 -1626
rect -2378 -1862 18986 -1626
rect 19222 -1862 54986 -1626
rect 55222 -1862 90986 -1626
rect 91222 -1862 126986 -1626
rect 127222 -1862 162986 -1626
rect 163222 -1862 198986 -1626
rect 199222 -1862 234986 -1626
rect 235222 -1862 270986 -1626
rect 271222 -1862 306986 -1626
rect 307222 -1862 342986 -1626
rect 343222 -1862 378986 -1626
rect 379222 -1862 414986 -1626
rect 415222 -1862 450986 -1626
rect 451222 -1862 486986 -1626
rect 487222 -1862 522986 -1626
rect 523222 -1862 558986 -1626
rect 559222 -1862 586302 -1626
rect 586538 -1862 586622 -1626
rect 586858 -1862 586890 -1626
rect -2966 -1894 586890 -1862
rect -3926 -2266 587850 -2234
rect -3926 -2502 -3894 -2266
rect -3658 -2502 -3574 -2266
rect -3338 -2502 4686 -2266
rect 4922 -2502 40686 -2266
rect 40922 -2502 76686 -2266
rect 76922 -2502 112686 -2266
rect 112922 -2502 148686 -2266
rect 148922 -2502 184686 -2266
rect 184922 -2502 220686 -2266
rect 220922 -2502 256686 -2266
rect 256922 -2502 292686 -2266
rect 292922 -2502 328686 -2266
rect 328922 -2502 364686 -2266
rect 364922 -2502 400686 -2266
rect 400922 -2502 436686 -2266
rect 436922 -2502 472686 -2266
rect 472922 -2502 508686 -2266
rect 508922 -2502 544686 -2266
rect 544922 -2502 580686 -2266
rect 580922 -2502 587262 -2266
rect 587498 -2502 587582 -2266
rect 587818 -2502 587850 -2266
rect -3926 -2586 587850 -2502
rect -3926 -2822 -3894 -2586
rect -3658 -2822 -3574 -2586
rect -3338 -2822 4686 -2586
rect 4922 -2822 40686 -2586
rect 40922 -2822 76686 -2586
rect 76922 -2822 112686 -2586
rect 112922 -2822 148686 -2586
rect 148922 -2822 184686 -2586
rect 184922 -2822 220686 -2586
rect 220922 -2822 256686 -2586
rect 256922 -2822 292686 -2586
rect 292922 -2822 328686 -2586
rect 328922 -2822 364686 -2586
rect 364922 -2822 400686 -2586
rect 400922 -2822 436686 -2586
rect 436922 -2822 472686 -2586
rect 472922 -2822 508686 -2586
rect 508922 -2822 544686 -2586
rect 544922 -2822 580686 -2586
rect 580922 -2822 587262 -2586
rect 587498 -2822 587582 -2586
rect 587818 -2822 587850 -2586
rect -3926 -2854 587850 -2822
rect -4886 -3226 588810 -3194
rect -4886 -3462 -4854 -3226
rect -4618 -3462 -4534 -3226
rect -4298 -3462 22686 -3226
rect 22922 -3462 58686 -3226
rect 58922 -3462 94686 -3226
rect 94922 -3462 130686 -3226
rect 130922 -3462 166686 -3226
rect 166922 -3462 202686 -3226
rect 202922 -3462 238686 -3226
rect 238922 -3462 274686 -3226
rect 274922 -3462 310686 -3226
rect 310922 -3462 346686 -3226
rect 346922 -3462 382686 -3226
rect 382922 -3462 418686 -3226
rect 418922 -3462 454686 -3226
rect 454922 -3462 490686 -3226
rect 490922 -3462 526686 -3226
rect 526922 -3462 562686 -3226
rect 562922 -3462 588222 -3226
rect 588458 -3462 588542 -3226
rect 588778 -3462 588810 -3226
rect -4886 -3546 588810 -3462
rect -4886 -3782 -4854 -3546
rect -4618 -3782 -4534 -3546
rect -4298 -3782 22686 -3546
rect 22922 -3782 58686 -3546
rect 58922 -3782 94686 -3546
rect 94922 -3782 130686 -3546
rect 130922 -3782 166686 -3546
rect 166922 -3782 202686 -3546
rect 202922 -3782 238686 -3546
rect 238922 -3782 274686 -3546
rect 274922 -3782 310686 -3546
rect 310922 -3782 346686 -3546
rect 346922 -3782 382686 -3546
rect 382922 -3782 418686 -3546
rect 418922 -3782 454686 -3546
rect 454922 -3782 490686 -3546
rect 490922 -3782 526686 -3546
rect 526922 -3782 562686 -3546
rect 562922 -3782 588222 -3546
rect 588458 -3782 588542 -3546
rect 588778 -3782 588810 -3546
rect -4886 -3814 588810 -3782
rect -5846 -4186 589770 -4154
rect -5846 -4422 -5814 -4186
rect -5578 -4422 -5494 -4186
rect -5258 -4422 8386 -4186
rect 8622 -4422 44386 -4186
rect 44622 -4422 80386 -4186
rect 80622 -4422 116386 -4186
rect 116622 -4422 152386 -4186
rect 152622 -4422 188386 -4186
rect 188622 -4422 224386 -4186
rect 224622 -4422 260386 -4186
rect 260622 -4422 296386 -4186
rect 296622 -4422 332386 -4186
rect 332622 -4422 368386 -4186
rect 368622 -4422 404386 -4186
rect 404622 -4422 440386 -4186
rect 440622 -4422 476386 -4186
rect 476622 -4422 512386 -4186
rect 512622 -4422 548386 -4186
rect 548622 -4422 589182 -4186
rect 589418 -4422 589502 -4186
rect 589738 -4422 589770 -4186
rect -5846 -4506 589770 -4422
rect -5846 -4742 -5814 -4506
rect -5578 -4742 -5494 -4506
rect -5258 -4742 8386 -4506
rect 8622 -4742 44386 -4506
rect 44622 -4742 80386 -4506
rect 80622 -4742 116386 -4506
rect 116622 -4742 152386 -4506
rect 152622 -4742 188386 -4506
rect 188622 -4742 224386 -4506
rect 224622 -4742 260386 -4506
rect 260622 -4742 296386 -4506
rect 296622 -4742 332386 -4506
rect 332622 -4742 368386 -4506
rect 368622 -4742 404386 -4506
rect 404622 -4742 440386 -4506
rect 440622 -4742 476386 -4506
rect 476622 -4742 512386 -4506
rect 512622 -4742 548386 -4506
rect 548622 -4742 589182 -4506
rect 589418 -4742 589502 -4506
rect 589738 -4742 589770 -4506
rect -5846 -4774 589770 -4742
rect -6806 -5146 590730 -5114
rect -6806 -5382 -6774 -5146
rect -6538 -5382 -6454 -5146
rect -6218 -5382 26386 -5146
rect 26622 -5382 62386 -5146
rect 62622 -5382 98386 -5146
rect 98622 -5382 134386 -5146
rect 134622 -5382 170386 -5146
rect 170622 -5382 206386 -5146
rect 206622 -5382 242386 -5146
rect 242622 -5382 278386 -5146
rect 278622 -5382 314386 -5146
rect 314622 -5382 350386 -5146
rect 350622 -5382 386386 -5146
rect 386622 -5382 422386 -5146
rect 422622 -5382 458386 -5146
rect 458622 -5382 494386 -5146
rect 494622 -5382 530386 -5146
rect 530622 -5382 566386 -5146
rect 566622 -5382 590142 -5146
rect 590378 -5382 590462 -5146
rect 590698 -5382 590730 -5146
rect -6806 -5466 590730 -5382
rect -6806 -5702 -6774 -5466
rect -6538 -5702 -6454 -5466
rect -6218 -5702 26386 -5466
rect 26622 -5702 62386 -5466
rect 62622 -5702 98386 -5466
rect 98622 -5702 134386 -5466
rect 134622 -5702 170386 -5466
rect 170622 -5702 206386 -5466
rect 206622 -5702 242386 -5466
rect 242622 -5702 278386 -5466
rect 278622 -5702 314386 -5466
rect 314622 -5702 350386 -5466
rect 350622 -5702 386386 -5466
rect 386622 -5702 422386 -5466
rect 422622 -5702 458386 -5466
rect 458622 -5702 494386 -5466
rect 494622 -5702 530386 -5466
rect 530622 -5702 566386 -5466
rect 566622 -5702 590142 -5466
rect 590378 -5702 590462 -5466
rect 590698 -5702 590730 -5466
rect -6806 -5734 590730 -5702
rect -7766 -6106 591690 -6074
rect -7766 -6342 -7734 -6106
rect -7498 -6342 -7414 -6106
rect -7178 -6342 12086 -6106
rect 12322 -6342 48086 -6106
rect 48322 -6342 84086 -6106
rect 84322 -6342 120086 -6106
rect 120322 -6342 156086 -6106
rect 156322 -6342 192086 -6106
rect 192322 -6342 228086 -6106
rect 228322 -6342 264086 -6106
rect 264322 -6342 300086 -6106
rect 300322 -6342 336086 -6106
rect 336322 -6342 372086 -6106
rect 372322 -6342 408086 -6106
rect 408322 -6342 444086 -6106
rect 444322 -6342 480086 -6106
rect 480322 -6342 516086 -6106
rect 516322 -6342 552086 -6106
rect 552322 -6342 591102 -6106
rect 591338 -6342 591422 -6106
rect 591658 -6342 591690 -6106
rect -7766 -6426 591690 -6342
rect -7766 -6662 -7734 -6426
rect -7498 -6662 -7414 -6426
rect -7178 -6662 12086 -6426
rect 12322 -6662 48086 -6426
rect 48322 -6662 84086 -6426
rect 84322 -6662 120086 -6426
rect 120322 -6662 156086 -6426
rect 156322 -6662 192086 -6426
rect 192322 -6662 228086 -6426
rect 228322 -6662 264086 -6426
rect 264322 -6662 300086 -6426
rect 300322 -6662 336086 -6426
rect 336322 -6662 372086 -6426
rect 372322 -6662 408086 -6426
rect 408322 -6662 444086 -6426
rect 444322 -6662 480086 -6426
rect 480322 -6662 516086 -6426
rect 516322 -6662 552086 -6426
rect 552322 -6662 591102 -6426
rect 591338 -6662 591422 -6426
rect 591658 -6662 591690 -6426
rect -7766 -6694 591690 -6662
rect -8726 -7066 592650 -7034
rect -8726 -7302 -8694 -7066
rect -8458 -7302 -8374 -7066
rect -8138 -7302 30086 -7066
rect 30322 -7302 66086 -7066
rect 66322 -7302 102086 -7066
rect 102322 -7302 138086 -7066
rect 138322 -7302 174086 -7066
rect 174322 -7302 210086 -7066
rect 210322 -7302 246086 -7066
rect 246322 -7302 282086 -7066
rect 282322 -7302 318086 -7066
rect 318322 -7302 354086 -7066
rect 354322 -7302 390086 -7066
rect 390322 -7302 426086 -7066
rect 426322 -7302 462086 -7066
rect 462322 -7302 498086 -7066
rect 498322 -7302 534086 -7066
rect 534322 -7302 570086 -7066
rect 570322 -7302 592062 -7066
rect 592298 -7302 592382 -7066
rect 592618 -7302 592650 -7066
rect -8726 -7386 592650 -7302
rect -8726 -7622 -8694 -7386
rect -8458 -7622 -8374 -7386
rect -8138 -7622 30086 -7386
rect 30322 -7622 66086 -7386
rect 66322 -7622 102086 -7386
rect 102322 -7622 138086 -7386
rect 138322 -7622 174086 -7386
rect 174322 -7622 210086 -7386
rect 210322 -7622 246086 -7386
rect 246322 -7622 282086 -7386
rect 282322 -7622 318086 -7386
rect 318322 -7622 354086 -7386
rect 354322 -7622 390086 -7386
rect 390322 -7622 426086 -7386
rect 426322 -7622 462086 -7386
rect 462322 -7622 498086 -7386
rect 498322 -7622 534086 -7386
rect 534322 -7622 570086 -7386
rect 570322 -7622 592062 -7386
rect 592298 -7622 592382 -7386
rect 592618 -7622 592650 -7386
rect -8726 -7654 592650 -7622
use sky130_sram_2kbyte_1rw1r_32x512_8  sram1
timestamp 1645590684
transform 1 0 340000 0 1 340000
box 0 0 136620 83308
use sky130_sram_2kbyte_1rw1r_32x512_8  sram
timestamp 1645590684
transform 1 0 40000 0 1 340000
box 0 0 136620 83308
use user_proj  mprj
timestamp 1645590684
transform 1 0 40000 0 1 40000
box 0 0 199424 201568
<< labels >>
rlabel metal3 s 583520 285276 584960 285516 6 analog_io[0]
port 0 nsew signal bidirectional
rlabel metal2 s 446098 703520 446210 704960 6 analog_io[10]
port 1 nsew signal bidirectional
rlabel metal2 s 381146 703520 381258 704960 6 analog_io[11]
port 2 nsew signal bidirectional
rlabel metal2 s 316286 703520 316398 704960 6 analog_io[12]
port 3 nsew signal bidirectional
rlabel metal2 s 251426 703520 251538 704960 6 analog_io[13]
port 4 nsew signal bidirectional
rlabel metal2 s 186474 703520 186586 704960 6 analog_io[14]
port 5 nsew signal bidirectional
rlabel metal2 s 121614 703520 121726 704960 6 analog_io[15]
port 6 nsew signal bidirectional
rlabel metal2 s 56754 703520 56866 704960 6 analog_io[16]
port 7 nsew signal bidirectional
rlabel metal3 s -960 697220 480 697460 4 analog_io[17]
port 8 nsew signal bidirectional
rlabel metal3 s -960 644996 480 645236 4 analog_io[18]
port 9 nsew signal bidirectional
rlabel metal3 s -960 592908 480 593148 4 analog_io[19]
port 10 nsew signal bidirectional
rlabel metal3 s 583520 338452 584960 338692 6 analog_io[1]
port 11 nsew signal bidirectional
rlabel metal3 s -960 540684 480 540924 4 analog_io[20]
port 12 nsew signal bidirectional
rlabel metal3 s -960 488596 480 488836 4 analog_io[21]
port 13 nsew signal bidirectional
rlabel metal3 s -960 436508 480 436748 4 analog_io[22]
port 14 nsew signal bidirectional
rlabel metal3 s -960 384284 480 384524 4 analog_io[23]
port 15 nsew signal bidirectional
rlabel metal3 s -960 332196 480 332436 4 analog_io[24]
port 16 nsew signal bidirectional
rlabel metal3 s -960 279972 480 280212 4 analog_io[25]
port 17 nsew signal bidirectional
rlabel metal3 s -960 227884 480 228124 4 analog_io[26]
port 18 nsew signal bidirectional
rlabel metal3 s -960 175796 480 176036 4 analog_io[27]
port 19 nsew signal bidirectional
rlabel metal3 s -960 123572 480 123812 4 analog_io[28]
port 20 nsew signal bidirectional
rlabel metal3 s 583520 391628 584960 391868 6 analog_io[2]
port 21 nsew signal bidirectional
rlabel metal3 s 583520 444668 584960 444908 6 analog_io[3]
port 22 nsew signal bidirectional
rlabel metal3 s 583520 497844 584960 498084 6 analog_io[4]
port 23 nsew signal bidirectional
rlabel metal3 s 583520 551020 584960 551260 6 analog_io[5]
port 24 nsew signal bidirectional
rlabel metal3 s 583520 604060 584960 604300 6 analog_io[6]
port 25 nsew signal bidirectional
rlabel metal3 s 583520 657236 584960 657476 6 analog_io[7]
port 26 nsew signal bidirectional
rlabel metal2 s 575818 703520 575930 704960 6 analog_io[8]
port 27 nsew signal bidirectional
rlabel metal2 s 510958 703520 511070 704960 6 analog_io[9]
port 28 nsew signal bidirectional
rlabel metal3 s 583520 6476 584960 6716 6 io_in[0]
port 29 nsew signal input
rlabel metal3 s 583520 457996 584960 458236 6 io_in[10]
port 30 nsew signal input
rlabel metal3 s 583520 511172 584960 511412 6 io_in[11]
port 31 nsew signal input
rlabel metal3 s 583520 564212 584960 564452 6 io_in[12]
port 32 nsew signal input
rlabel metal3 s 583520 617388 584960 617628 6 io_in[13]
port 33 nsew signal input
rlabel metal3 s 583520 670564 584960 670804 6 io_in[14]
port 34 nsew signal input
rlabel metal2 s 559626 703520 559738 704960 6 io_in[15]
port 35 nsew signal input
rlabel metal2 s 494766 703520 494878 704960 6 io_in[16]
port 36 nsew signal input
rlabel metal2 s 429814 703520 429926 704960 6 io_in[17]
port 37 nsew signal input
rlabel metal2 s 364954 703520 365066 704960 6 io_in[18]
port 38 nsew signal input
rlabel metal2 s 300094 703520 300206 704960 6 io_in[19]
port 39 nsew signal input
rlabel metal3 s 583520 46188 584960 46428 6 io_in[1]
port 40 nsew signal input
rlabel metal2 s 235142 703520 235254 704960 6 io_in[20]
port 41 nsew signal input
rlabel metal2 s 170282 703520 170394 704960 6 io_in[21]
port 42 nsew signal input
rlabel metal2 s 105422 703520 105534 704960 6 io_in[22]
port 43 nsew signal input
rlabel metal2 s 40470 703520 40582 704960 6 io_in[23]
port 44 nsew signal input
rlabel metal3 s -960 684164 480 684404 4 io_in[24]
port 45 nsew signal input
rlabel metal3 s -960 631940 480 632180 4 io_in[25]
port 46 nsew signal input
rlabel metal3 s -960 579852 480 580092 4 io_in[26]
port 47 nsew signal input
rlabel metal3 s -960 527764 480 528004 4 io_in[27]
port 48 nsew signal input
rlabel metal3 s -960 475540 480 475780 4 io_in[28]
port 49 nsew signal input
rlabel metal3 s -960 423452 480 423692 4 io_in[29]
port 50 nsew signal input
rlabel metal3 s 583520 86036 584960 86276 6 io_in[2]
port 51 nsew signal input
rlabel metal3 s -960 371228 480 371468 4 io_in[30]
port 52 nsew signal input
rlabel metal3 s -960 319140 480 319380 4 io_in[31]
port 53 nsew signal input
rlabel metal3 s -960 267052 480 267292 4 io_in[32]
port 54 nsew signal input
rlabel metal3 s -960 214828 480 215068 4 io_in[33]
port 55 nsew signal input
rlabel metal3 s -960 162740 480 162980 4 io_in[34]
port 56 nsew signal input
rlabel metal3 s -960 110516 480 110756 4 io_in[35]
port 57 nsew signal input
rlabel metal3 s -960 71484 480 71724 4 io_in[36]
port 58 nsew signal input
rlabel metal3 s -960 32316 480 32556 4 io_in[37]
port 59 nsew signal input
rlabel metal3 s 583520 125884 584960 126124 6 io_in[3]
port 60 nsew signal input
rlabel metal3 s 583520 165732 584960 165972 6 io_in[4]
port 61 nsew signal input
rlabel metal3 s 583520 205580 584960 205820 6 io_in[5]
port 62 nsew signal input
rlabel metal3 s 583520 245428 584960 245668 6 io_in[6]
port 63 nsew signal input
rlabel metal3 s 583520 298604 584960 298844 6 io_in[7]
port 64 nsew signal input
rlabel metal3 s 583520 351780 584960 352020 6 io_in[8]
port 65 nsew signal input
rlabel metal3 s 583520 404820 584960 405060 6 io_in[9]
port 66 nsew signal input
rlabel metal3 s 583520 32996 584960 33236 6 io_oeb[0]
port 67 nsew signal tristate
rlabel metal3 s 583520 484516 584960 484756 6 io_oeb[10]
port 68 nsew signal tristate
rlabel metal3 s 583520 537692 584960 537932 6 io_oeb[11]
port 69 nsew signal tristate
rlabel metal3 s 583520 590868 584960 591108 6 io_oeb[12]
port 70 nsew signal tristate
rlabel metal3 s 583520 643908 584960 644148 6 io_oeb[13]
port 71 nsew signal tristate
rlabel metal3 s 583520 697084 584960 697324 6 io_oeb[14]
port 72 nsew signal tristate
rlabel metal2 s 527150 703520 527262 704960 6 io_oeb[15]
port 73 nsew signal tristate
rlabel metal2 s 462290 703520 462402 704960 6 io_oeb[16]
port 74 nsew signal tristate
rlabel metal2 s 397430 703520 397542 704960 6 io_oeb[17]
port 75 nsew signal tristate
rlabel metal2 s 332478 703520 332590 704960 6 io_oeb[18]
port 76 nsew signal tristate
rlabel metal2 s 267618 703520 267730 704960 6 io_oeb[19]
port 77 nsew signal tristate
rlabel metal3 s 583520 72844 584960 73084 6 io_oeb[1]
port 78 nsew signal tristate
rlabel metal2 s 202758 703520 202870 704960 6 io_oeb[20]
port 79 nsew signal tristate
rlabel metal2 s 137806 703520 137918 704960 6 io_oeb[21]
port 80 nsew signal tristate
rlabel metal2 s 72946 703520 73058 704960 6 io_oeb[22]
port 81 nsew signal tristate
rlabel metal2 s 8086 703520 8198 704960 6 io_oeb[23]
port 82 nsew signal tristate
rlabel metal3 s -960 658052 480 658292 4 io_oeb[24]
port 83 nsew signal tristate
rlabel metal3 s -960 605964 480 606204 4 io_oeb[25]
port 84 nsew signal tristate
rlabel metal3 s -960 553740 480 553980 4 io_oeb[26]
port 85 nsew signal tristate
rlabel metal3 s -960 501652 480 501892 4 io_oeb[27]
port 86 nsew signal tristate
rlabel metal3 s -960 449428 480 449668 4 io_oeb[28]
port 87 nsew signal tristate
rlabel metal3 s -960 397340 480 397580 4 io_oeb[29]
port 88 nsew signal tristate
rlabel metal3 s 583520 112692 584960 112932 6 io_oeb[2]
port 89 nsew signal tristate
rlabel metal3 s -960 345252 480 345492 4 io_oeb[30]
port 90 nsew signal tristate
rlabel metal3 s -960 293028 480 293268 4 io_oeb[31]
port 91 nsew signal tristate
rlabel metal3 s -960 240940 480 241180 4 io_oeb[32]
port 92 nsew signal tristate
rlabel metal3 s -960 188716 480 188956 4 io_oeb[33]
port 93 nsew signal tristate
rlabel metal3 s -960 136628 480 136868 4 io_oeb[34]
port 94 nsew signal tristate
rlabel metal3 s -960 84540 480 84780 4 io_oeb[35]
port 95 nsew signal tristate
rlabel metal3 s -960 45372 480 45612 4 io_oeb[36]
port 96 nsew signal tristate
rlabel metal3 s -960 6340 480 6580 4 io_oeb[37]
port 97 nsew signal tristate
rlabel metal3 s 583520 152540 584960 152780 6 io_oeb[3]
port 98 nsew signal tristate
rlabel metal3 s 583520 192388 584960 192628 6 io_oeb[4]
port 99 nsew signal tristate
rlabel metal3 s 583520 232236 584960 232476 6 io_oeb[5]
port 100 nsew signal tristate
rlabel metal3 s 583520 272084 584960 272324 6 io_oeb[6]
port 101 nsew signal tristate
rlabel metal3 s 583520 325124 584960 325364 6 io_oeb[7]
port 102 nsew signal tristate
rlabel metal3 s 583520 378300 584960 378540 6 io_oeb[8]
port 103 nsew signal tristate
rlabel metal3 s 583520 431476 584960 431716 6 io_oeb[9]
port 104 nsew signal tristate
rlabel metal3 s 583520 19668 584960 19908 6 io_out[0]
port 105 nsew signal tristate
rlabel metal3 s 583520 471324 584960 471564 6 io_out[10]
port 106 nsew signal tristate
rlabel metal3 s 583520 524364 584960 524604 6 io_out[11]
port 107 nsew signal tristate
rlabel metal3 s 583520 577540 584960 577780 6 io_out[12]
port 108 nsew signal tristate
rlabel metal3 s 583520 630716 584960 630956 6 io_out[13]
port 109 nsew signal tristate
rlabel metal3 s 583520 683756 584960 683996 6 io_out[14]
port 110 nsew signal tristate
rlabel metal2 s 543434 703520 543546 704960 6 io_out[15]
port 111 nsew signal tristate
rlabel metal2 s 478482 703520 478594 704960 6 io_out[16]
port 112 nsew signal tristate
rlabel metal2 s 413622 703520 413734 704960 6 io_out[17]
port 113 nsew signal tristate
rlabel metal2 s 348762 703520 348874 704960 6 io_out[18]
port 114 nsew signal tristate
rlabel metal2 s 283810 703520 283922 704960 6 io_out[19]
port 115 nsew signal tristate
rlabel metal3 s 583520 59516 584960 59756 6 io_out[1]
port 116 nsew signal tristate
rlabel metal2 s 218950 703520 219062 704960 6 io_out[20]
port 117 nsew signal tristate
rlabel metal2 s 154090 703520 154202 704960 6 io_out[21]
port 118 nsew signal tristate
rlabel metal2 s 89138 703520 89250 704960 6 io_out[22]
port 119 nsew signal tristate
rlabel metal2 s 24278 703520 24390 704960 6 io_out[23]
port 120 nsew signal tristate
rlabel metal3 s -960 671108 480 671348 4 io_out[24]
port 121 nsew signal tristate
rlabel metal3 s -960 619020 480 619260 4 io_out[25]
port 122 nsew signal tristate
rlabel metal3 s -960 566796 480 567036 4 io_out[26]
port 123 nsew signal tristate
rlabel metal3 s -960 514708 480 514948 4 io_out[27]
port 124 nsew signal tristate
rlabel metal3 s -960 462484 480 462724 4 io_out[28]
port 125 nsew signal tristate
rlabel metal3 s -960 410396 480 410636 4 io_out[29]
port 126 nsew signal tristate
rlabel metal3 s 583520 99364 584960 99604 6 io_out[2]
port 127 nsew signal tristate
rlabel metal3 s -960 358308 480 358548 4 io_out[30]
port 128 nsew signal tristate
rlabel metal3 s -960 306084 480 306324 4 io_out[31]
port 129 nsew signal tristate
rlabel metal3 s -960 253996 480 254236 4 io_out[32]
port 130 nsew signal tristate
rlabel metal3 s -960 201772 480 202012 4 io_out[33]
port 131 nsew signal tristate
rlabel metal3 s -960 149684 480 149924 4 io_out[34]
port 132 nsew signal tristate
rlabel metal3 s -960 97460 480 97700 4 io_out[35]
port 133 nsew signal tristate
rlabel metal3 s -960 58428 480 58668 4 io_out[36]
port 134 nsew signal tristate
rlabel metal3 s -960 19260 480 19500 4 io_out[37]
port 135 nsew signal tristate
rlabel metal3 s 583520 139212 584960 139452 6 io_out[3]
port 136 nsew signal tristate
rlabel metal3 s 583520 179060 584960 179300 6 io_out[4]
port 137 nsew signal tristate
rlabel metal3 s 583520 218908 584960 219148 6 io_out[5]
port 138 nsew signal tristate
rlabel metal3 s 583520 258756 584960 258996 6 io_out[6]
port 139 nsew signal tristate
rlabel metal3 s 583520 311932 584960 312172 6 io_out[7]
port 140 nsew signal tristate
rlabel metal3 s 583520 364972 584960 365212 6 io_out[8]
port 141 nsew signal tristate
rlabel metal3 s 583520 418148 584960 418388 6 io_out[9]
port 142 nsew signal tristate
rlabel metal2 s 125846 -960 125958 480 8 la_data_in[0]
port 143 nsew signal input
rlabel metal2 s 480506 -960 480618 480 8 la_data_in[100]
port 144 nsew signal input
rlabel metal2 s 484002 -960 484114 480 8 la_data_in[101]
port 145 nsew signal input
rlabel metal2 s 487590 -960 487702 480 8 la_data_in[102]
port 146 nsew signal input
rlabel metal2 s 491086 -960 491198 480 8 la_data_in[103]
port 147 nsew signal input
rlabel metal2 s 494674 -960 494786 480 8 la_data_in[104]
port 148 nsew signal input
rlabel metal2 s 498170 -960 498282 480 8 la_data_in[105]
port 149 nsew signal input
rlabel metal2 s 501758 -960 501870 480 8 la_data_in[106]
port 150 nsew signal input
rlabel metal2 s 505346 -960 505458 480 8 la_data_in[107]
port 151 nsew signal input
rlabel metal2 s 508842 -960 508954 480 8 la_data_in[108]
port 152 nsew signal input
rlabel metal2 s 512430 -960 512542 480 8 la_data_in[109]
port 153 nsew signal input
rlabel metal2 s 161266 -960 161378 480 8 la_data_in[10]
port 154 nsew signal input
rlabel metal2 s 515926 -960 516038 480 8 la_data_in[110]
port 155 nsew signal input
rlabel metal2 s 519514 -960 519626 480 8 la_data_in[111]
port 156 nsew signal input
rlabel metal2 s 523010 -960 523122 480 8 la_data_in[112]
port 157 nsew signal input
rlabel metal2 s 526598 -960 526710 480 8 la_data_in[113]
port 158 nsew signal input
rlabel metal2 s 530094 -960 530206 480 8 la_data_in[114]
port 159 nsew signal input
rlabel metal2 s 533682 -960 533794 480 8 la_data_in[115]
port 160 nsew signal input
rlabel metal2 s 537178 -960 537290 480 8 la_data_in[116]
port 161 nsew signal input
rlabel metal2 s 540766 -960 540878 480 8 la_data_in[117]
port 162 nsew signal input
rlabel metal2 s 544354 -960 544466 480 8 la_data_in[118]
port 163 nsew signal input
rlabel metal2 s 547850 -960 547962 480 8 la_data_in[119]
port 164 nsew signal input
rlabel metal2 s 164854 -960 164966 480 8 la_data_in[11]
port 165 nsew signal input
rlabel metal2 s 551438 -960 551550 480 8 la_data_in[120]
port 166 nsew signal input
rlabel metal2 s 554934 -960 555046 480 8 la_data_in[121]
port 167 nsew signal input
rlabel metal2 s 558522 -960 558634 480 8 la_data_in[122]
port 168 nsew signal input
rlabel metal2 s 562018 -960 562130 480 8 la_data_in[123]
port 169 nsew signal input
rlabel metal2 s 565606 -960 565718 480 8 la_data_in[124]
port 170 nsew signal input
rlabel metal2 s 569102 -960 569214 480 8 la_data_in[125]
port 171 nsew signal input
rlabel metal2 s 572690 -960 572802 480 8 la_data_in[126]
port 172 nsew signal input
rlabel metal2 s 576278 -960 576390 480 8 la_data_in[127]
port 173 nsew signal input
rlabel metal2 s 168350 -960 168462 480 8 la_data_in[12]
port 174 nsew signal input
rlabel metal2 s 171938 -960 172050 480 8 la_data_in[13]
port 175 nsew signal input
rlabel metal2 s 175434 -960 175546 480 8 la_data_in[14]
port 176 nsew signal input
rlabel metal2 s 179022 -960 179134 480 8 la_data_in[15]
port 177 nsew signal input
rlabel metal2 s 182518 -960 182630 480 8 la_data_in[16]
port 178 nsew signal input
rlabel metal2 s 186106 -960 186218 480 8 la_data_in[17]
port 179 nsew signal input
rlabel metal2 s 189694 -960 189806 480 8 la_data_in[18]
port 180 nsew signal input
rlabel metal2 s 193190 -960 193302 480 8 la_data_in[19]
port 181 nsew signal input
rlabel metal2 s 129342 -960 129454 480 8 la_data_in[1]
port 182 nsew signal input
rlabel metal2 s 196778 -960 196890 480 8 la_data_in[20]
port 183 nsew signal input
rlabel metal2 s 200274 -960 200386 480 8 la_data_in[21]
port 184 nsew signal input
rlabel metal2 s 203862 -960 203974 480 8 la_data_in[22]
port 185 nsew signal input
rlabel metal2 s 207358 -960 207470 480 8 la_data_in[23]
port 186 nsew signal input
rlabel metal2 s 210946 -960 211058 480 8 la_data_in[24]
port 187 nsew signal input
rlabel metal2 s 214442 -960 214554 480 8 la_data_in[25]
port 188 nsew signal input
rlabel metal2 s 218030 -960 218142 480 8 la_data_in[26]
port 189 nsew signal input
rlabel metal2 s 221526 -960 221638 480 8 la_data_in[27]
port 190 nsew signal input
rlabel metal2 s 225114 -960 225226 480 8 la_data_in[28]
port 191 nsew signal input
rlabel metal2 s 228702 -960 228814 480 8 la_data_in[29]
port 192 nsew signal input
rlabel metal2 s 132930 -960 133042 480 8 la_data_in[2]
port 193 nsew signal input
rlabel metal2 s 232198 -960 232310 480 8 la_data_in[30]
port 194 nsew signal input
rlabel metal2 s 235786 -960 235898 480 8 la_data_in[31]
port 195 nsew signal input
rlabel metal2 s 239282 -960 239394 480 8 la_data_in[32]
port 196 nsew signal input
rlabel metal2 s 242870 -960 242982 480 8 la_data_in[33]
port 197 nsew signal input
rlabel metal2 s 246366 -960 246478 480 8 la_data_in[34]
port 198 nsew signal input
rlabel metal2 s 249954 -960 250066 480 8 la_data_in[35]
port 199 nsew signal input
rlabel metal2 s 253450 -960 253562 480 8 la_data_in[36]
port 200 nsew signal input
rlabel metal2 s 257038 -960 257150 480 8 la_data_in[37]
port 201 nsew signal input
rlabel metal2 s 260626 -960 260738 480 8 la_data_in[38]
port 202 nsew signal input
rlabel metal2 s 264122 -960 264234 480 8 la_data_in[39]
port 203 nsew signal input
rlabel metal2 s 136426 -960 136538 480 8 la_data_in[3]
port 204 nsew signal input
rlabel metal2 s 267710 -960 267822 480 8 la_data_in[40]
port 205 nsew signal input
rlabel metal2 s 271206 -960 271318 480 8 la_data_in[41]
port 206 nsew signal input
rlabel metal2 s 274794 -960 274906 480 8 la_data_in[42]
port 207 nsew signal input
rlabel metal2 s 278290 -960 278402 480 8 la_data_in[43]
port 208 nsew signal input
rlabel metal2 s 281878 -960 281990 480 8 la_data_in[44]
port 209 nsew signal input
rlabel metal2 s 285374 -960 285486 480 8 la_data_in[45]
port 210 nsew signal input
rlabel metal2 s 288962 -960 289074 480 8 la_data_in[46]
port 211 nsew signal input
rlabel metal2 s 292550 -960 292662 480 8 la_data_in[47]
port 212 nsew signal input
rlabel metal2 s 296046 -960 296158 480 8 la_data_in[48]
port 213 nsew signal input
rlabel metal2 s 299634 -960 299746 480 8 la_data_in[49]
port 214 nsew signal input
rlabel metal2 s 140014 -960 140126 480 8 la_data_in[4]
port 215 nsew signal input
rlabel metal2 s 303130 -960 303242 480 8 la_data_in[50]
port 216 nsew signal input
rlabel metal2 s 306718 -960 306830 480 8 la_data_in[51]
port 217 nsew signal input
rlabel metal2 s 310214 -960 310326 480 8 la_data_in[52]
port 218 nsew signal input
rlabel metal2 s 313802 -960 313914 480 8 la_data_in[53]
port 219 nsew signal input
rlabel metal2 s 317298 -960 317410 480 8 la_data_in[54]
port 220 nsew signal input
rlabel metal2 s 320886 -960 320998 480 8 la_data_in[55]
port 221 nsew signal input
rlabel metal2 s 324382 -960 324494 480 8 la_data_in[56]
port 222 nsew signal input
rlabel metal2 s 327970 -960 328082 480 8 la_data_in[57]
port 223 nsew signal input
rlabel metal2 s 331558 -960 331670 480 8 la_data_in[58]
port 224 nsew signal input
rlabel metal2 s 335054 -960 335166 480 8 la_data_in[59]
port 225 nsew signal input
rlabel metal2 s 143510 -960 143622 480 8 la_data_in[5]
port 226 nsew signal input
rlabel metal2 s 338642 -960 338754 480 8 la_data_in[60]
port 227 nsew signal input
rlabel metal2 s 342138 -960 342250 480 8 la_data_in[61]
port 228 nsew signal input
rlabel metal2 s 345726 -960 345838 480 8 la_data_in[62]
port 229 nsew signal input
rlabel metal2 s 349222 -960 349334 480 8 la_data_in[63]
port 230 nsew signal input
rlabel metal2 s 352810 -960 352922 480 8 la_data_in[64]
port 231 nsew signal input
rlabel metal2 s 356306 -960 356418 480 8 la_data_in[65]
port 232 nsew signal input
rlabel metal2 s 359894 -960 360006 480 8 la_data_in[66]
port 233 nsew signal input
rlabel metal2 s 363482 -960 363594 480 8 la_data_in[67]
port 234 nsew signal input
rlabel metal2 s 366978 -960 367090 480 8 la_data_in[68]
port 235 nsew signal input
rlabel metal2 s 370566 -960 370678 480 8 la_data_in[69]
port 236 nsew signal input
rlabel metal2 s 147098 -960 147210 480 8 la_data_in[6]
port 237 nsew signal input
rlabel metal2 s 374062 -960 374174 480 8 la_data_in[70]
port 238 nsew signal input
rlabel metal2 s 377650 -960 377762 480 8 la_data_in[71]
port 239 nsew signal input
rlabel metal2 s 381146 -960 381258 480 8 la_data_in[72]
port 240 nsew signal input
rlabel metal2 s 384734 -960 384846 480 8 la_data_in[73]
port 241 nsew signal input
rlabel metal2 s 388230 -960 388342 480 8 la_data_in[74]
port 242 nsew signal input
rlabel metal2 s 391818 -960 391930 480 8 la_data_in[75]
port 243 nsew signal input
rlabel metal2 s 395314 -960 395426 480 8 la_data_in[76]
port 244 nsew signal input
rlabel metal2 s 398902 -960 399014 480 8 la_data_in[77]
port 245 nsew signal input
rlabel metal2 s 402490 -960 402602 480 8 la_data_in[78]
port 246 nsew signal input
rlabel metal2 s 405986 -960 406098 480 8 la_data_in[79]
port 247 nsew signal input
rlabel metal2 s 150594 -960 150706 480 8 la_data_in[7]
port 248 nsew signal input
rlabel metal2 s 409574 -960 409686 480 8 la_data_in[80]
port 249 nsew signal input
rlabel metal2 s 413070 -960 413182 480 8 la_data_in[81]
port 250 nsew signal input
rlabel metal2 s 416658 -960 416770 480 8 la_data_in[82]
port 251 nsew signal input
rlabel metal2 s 420154 -960 420266 480 8 la_data_in[83]
port 252 nsew signal input
rlabel metal2 s 423742 -960 423854 480 8 la_data_in[84]
port 253 nsew signal input
rlabel metal2 s 427238 -960 427350 480 8 la_data_in[85]
port 254 nsew signal input
rlabel metal2 s 430826 -960 430938 480 8 la_data_in[86]
port 255 nsew signal input
rlabel metal2 s 434414 -960 434526 480 8 la_data_in[87]
port 256 nsew signal input
rlabel metal2 s 437910 -960 438022 480 8 la_data_in[88]
port 257 nsew signal input
rlabel metal2 s 441498 -960 441610 480 8 la_data_in[89]
port 258 nsew signal input
rlabel metal2 s 154182 -960 154294 480 8 la_data_in[8]
port 259 nsew signal input
rlabel metal2 s 444994 -960 445106 480 8 la_data_in[90]
port 260 nsew signal input
rlabel metal2 s 448582 -960 448694 480 8 la_data_in[91]
port 261 nsew signal input
rlabel metal2 s 452078 -960 452190 480 8 la_data_in[92]
port 262 nsew signal input
rlabel metal2 s 455666 -960 455778 480 8 la_data_in[93]
port 263 nsew signal input
rlabel metal2 s 459162 -960 459274 480 8 la_data_in[94]
port 264 nsew signal input
rlabel metal2 s 462750 -960 462862 480 8 la_data_in[95]
port 265 nsew signal input
rlabel metal2 s 466246 -960 466358 480 8 la_data_in[96]
port 266 nsew signal input
rlabel metal2 s 469834 -960 469946 480 8 la_data_in[97]
port 267 nsew signal input
rlabel metal2 s 473422 -960 473534 480 8 la_data_in[98]
port 268 nsew signal input
rlabel metal2 s 476918 -960 477030 480 8 la_data_in[99]
port 269 nsew signal input
rlabel metal2 s 157770 -960 157882 480 8 la_data_in[9]
port 270 nsew signal input
rlabel metal2 s 126950 -960 127062 480 8 la_data_out[0]
port 271 nsew signal tristate
rlabel metal2 s 481702 -960 481814 480 8 la_data_out[100]
port 272 nsew signal tristate
rlabel metal2 s 485198 -960 485310 480 8 la_data_out[101]
port 273 nsew signal tristate
rlabel metal2 s 488786 -960 488898 480 8 la_data_out[102]
port 274 nsew signal tristate
rlabel metal2 s 492282 -960 492394 480 8 la_data_out[103]
port 275 nsew signal tristate
rlabel metal2 s 495870 -960 495982 480 8 la_data_out[104]
port 276 nsew signal tristate
rlabel metal2 s 499366 -960 499478 480 8 la_data_out[105]
port 277 nsew signal tristate
rlabel metal2 s 502954 -960 503066 480 8 la_data_out[106]
port 278 nsew signal tristate
rlabel metal2 s 506450 -960 506562 480 8 la_data_out[107]
port 279 nsew signal tristate
rlabel metal2 s 510038 -960 510150 480 8 la_data_out[108]
port 280 nsew signal tristate
rlabel metal2 s 513534 -960 513646 480 8 la_data_out[109]
port 281 nsew signal tristate
rlabel metal2 s 162462 -960 162574 480 8 la_data_out[10]
port 282 nsew signal tristate
rlabel metal2 s 517122 -960 517234 480 8 la_data_out[110]
port 283 nsew signal tristate
rlabel metal2 s 520710 -960 520822 480 8 la_data_out[111]
port 284 nsew signal tristate
rlabel metal2 s 524206 -960 524318 480 8 la_data_out[112]
port 285 nsew signal tristate
rlabel metal2 s 527794 -960 527906 480 8 la_data_out[113]
port 286 nsew signal tristate
rlabel metal2 s 531290 -960 531402 480 8 la_data_out[114]
port 287 nsew signal tristate
rlabel metal2 s 534878 -960 534990 480 8 la_data_out[115]
port 288 nsew signal tristate
rlabel metal2 s 538374 -960 538486 480 8 la_data_out[116]
port 289 nsew signal tristate
rlabel metal2 s 541962 -960 542074 480 8 la_data_out[117]
port 290 nsew signal tristate
rlabel metal2 s 545458 -960 545570 480 8 la_data_out[118]
port 291 nsew signal tristate
rlabel metal2 s 549046 -960 549158 480 8 la_data_out[119]
port 292 nsew signal tristate
rlabel metal2 s 166050 -960 166162 480 8 la_data_out[11]
port 293 nsew signal tristate
rlabel metal2 s 552634 -960 552746 480 8 la_data_out[120]
port 294 nsew signal tristate
rlabel metal2 s 556130 -960 556242 480 8 la_data_out[121]
port 295 nsew signal tristate
rlabel metal2 s 559718 -960 559830 480 8 la_data_out[122]
port 296 nsew signal tristate
rlabel metal2 s 563214 -960 563326 480 8 la_data_out[123]
port 297 nsew signal tristate
rlabel metal2 s 566802 -960 566914 480 8 la_data_out[124]
port 298 nsew signal tristate
rlabel metal2 s 570298 -960 570410 480 8 la_data_out[125]
port 299 nsew signal tristate
rlabel metal2 s 573886 -960 573998 480 8 la_data_out[126]
port 300 nsew signal tristate
rlabel metal2 s 577382 -960 577494 480 8 la_data_out[127]
port 301 nsew signal tristate
rlabel metal2 s 169546 -960 169658 480 8 la_data_out[12]
port 302 nsew signal tristate
rlabel metal2 s 173134 -960 173246 480 8 la_data_out[13]
port 303 nsew signal tristate
rlabel metal2 s 176630 -960 176742 480 8 la_data_out[14]
port 304 nsew signal tristate
rlabel metal2 s 180218 -960 180330 480 8 la_data_out[15]
port 305 nsew signal tristate
rlabel metal2 s 183714 -960 183826 480 8 la_data_out[16]
port 306 nsew signal tristate
rlabel metal2 s 187302 -960 187414 480 8 la_data_out[17]
port 307 nsew signal tristate
rlabel metal2 s 190798 -960 190910 480 8 la_data_out[18]
port 308 nsew signal tristate
rlabel metal2 s 194386 -960 194498 480 8 la_data_out[19]
port 309 nsew signal tristate
rlabel metal2 s 130538 -960 130650 480 8 la_data_out[1]
port 310 nsew signal tristate
rlabel metal2 s 197882 -960 197994 480 8 la_data_out[20]
port 311 nsew signal tristate
rlabel metal2 s 201470 -960 201582 480 8 la_data_out[21]
port 312 nsew signal tristate
rlabel metal2 s 205058 -960 205170 480 8 la_data_out[22]
port 313 nsew signal tristate
rlabel metal2 s 208554 -960 208666 480 8 la_data_out[23]
port 314 nsew signal tristate
rlabel metal2 s 212142 -960 212254 480 8 la_data_out[24]
port 315 nsew signal tristate
rlabel metal2 s 215638 -960 215750 480 8 la_data_out[25]
port 316 nsew signal tristate
rlabel metal2 s 219226 -960 219338 480 8 la_data_out[26]
port 317 nsew signal tristate
rlabel metal2 s 222722 -960 222834 480 8 la_data_out[27]
port 318 nsew signal tristate
rlabel metal2 s 226310 -960 226422 480 8 la_data_out[28]
port 319 nsew signal tristate
rlabel metal2 s 229806 -960 229918 480 8 la_data_out[29]
port 320 nsew signal tristate
rlabel metal2 s 134126 -960 134238 480 8 la_data_out[2]
port 321 nsew signal tristate
rlabel metal2 s 233394 -960 233506 480 8 la_data_out[30]
port 322 nsew signal tristate
rlabel metal2 s 236982 -960 237094 480 8 la_data_out[31]
port 323 nsew signal tristate
rlabel metal2 s 240478 -960 240590 480 8 la_data_out[32]
port 324 nsew signal tristate
rlabel metal2 s 244066 -960 244178 480 8 la_data_out[33]
port 325 nsew signal tristate
rlabel metal2 s 247562 -960 247674 480 8 la_data_out[34]
port 326 nsew signal tristate
rlabel metal2 s 251150 -960 251262 480 8 la_data_out[35]
port 327 nsew signal tristate
rlabel metal2 s 254646 -960 254758 480 8 la_data_out[36]
port 328 nsew signal tristate
rlabel metal2 s 258234 -960 258346 480 8 la_data_out[37]
port 329 nsew signal tristate
rlabel metal2 s 261730 -960 261842 480 8 la_data_out[38]
port 330 nsew signal tristate
rlabel metal2 s 265318 -960 265430 480 8 la_data_out[39]
port 331 nsew signal tristate
rlabel metal2 s 137622 -960 137734 480 8 la_data_out[3]
port 332 nsew signal tristate
rlabel metal2 s 268814 -960 268926 480 8 la_data_out[40]
port 333 nsew signal tristate
rlabel metal2 s 272402 -960 272514 480 8 la_data_out[41]
port 334 nsew signal tristate
rlabel metal2 s 275990 -960 276102 480 8 la_data_out[42]
port 335 nsew signal tristate
rlabel metal2 s 279486 -960 279598 480 8 la_data_out[43]
port 336 nsew signal tristate
rlabel metal2 s 283074 -960 283186 480 8 la_data_out[44]
port 337 nsew signal tristate
rlabel metal2 s 286570 -960 286682 480 8 la_data_out[45]
port 338 nsew signal tristate
rlabel metal2 s 290158 -960 290270 480 8 la_data_out[46]
port 339 nsew signal tristate
rlabel metal2 s 293654 -960 293766 480 8 la_data_out[47]
port 340 nsew signal tristate
rlabel metal2 s 297242 -960 297354 480 8 la_data_out[48]
port 341 nsew signal tristate
rlabel metal2 s 300738 -960 300850 480 8 la_data_out[49]
port 342 nsew signal tristate
rlabel metal2 s 141210 -960 141322 480 8 la_data_out[4]
port 343 nsew signal tristate
rlabel metal2 s 304326 -960 304438 480 8 la_data_out[50]
port 344 nsew signal tristate
rlabel metal2 s 307914 -960 308026 480 8 la_data_out[51]
port 345 nsew signal tristate
rlabel metal2 s 311410 -960 311522 480 8 la_data_out[52]
port 346 nsew signal tristate
rlabel metal2 s 314998 -960 315110 480 8 la_data_out[53]
port 347 nsew signal tristate
rlabel metal2 s 318494 -960 318606 480 8 la_data_out[54]
port 348 nsew signal tristate
rlabel metal2 s 322082 -960 322194 480 8 la_data_out[55]
port 349 nsew signal tristate
rlabel metal2 s 325578 -960 325690 480 8 la_data_out[56]
port 350 nsew signal tristate
rlabel metal2 s 329166 -960 329278 480 8 la_data_out[57]
port 351 nsew signal tristate
rlabel metal2 s 332662 -960 332774 480 8 la_data_out[58]
port 352 nsew signal tristate
rlabel metal2 s 336250 -960 336362 480 8 la_data_out[59]
port 353 nsew signal tristate
rlabel metal2 s 144706 -960 144818 480 8 la_data_out[5]
port 354 nsew signal tristate
rlabel metal2 s 339838 -960 339950 480 8 la_data_out[60]
port 355 nsew signal tristate
rlabel metal2 s 343334 -960 343446 480 8 la_data_out[61]
port 356 nsew signal tristate
rlabel metal2 s 346922 -960 347034 480 8 la_data_out[62]
port 357 nsew signal tristate
rlabel metal2 s 350418 -960 350530 480 8 la_data_out[63]
port 358 nsew signal tristate
rlabel metal2 s 354006 -960 354118 480 8 la_data_out[64]
port 359 nsew signal tristate
rlabel metal2 s 357502 -960 357614 480 8 la_data_out[65]
port 360 nsew signal tristate
rlabel metal2 s 361090 -960 361202 480 8 la_data_out[66]
port 361 nsew signal tristate
rlabel metal2 s 364586 -960 364698 480 8 la_data_out[67]
port 362 nsew signal tristate
rlabel metal2 s 368174 -960 368286 480 8 la_data_out[68]
port 363 nsew signal tristate
rlabel metal2 s 371670 -960 371782 480 8 la_data_out[69]
port 364 nsew signal tristate
rlabel metal2 s 148294 -960 148406 480 8 la_data_out[6]
port 365 nsew signal tristate
rlabel metal2 s 375258 -960 375370 480 8 la_data_out[70]
port 366 nsew signal tristate
rlabel metal2 s 378846 -960 378958 480 8 la_data_out[71]
port 367 nsew signal tristate
rlabel metal2 s 382342 -960 382454 480 8 la_data_out[72]
port 368 nsew signal tristate
rlabel metal2 s 385930 -960 386042 480 8 la_data_out[73]
port 369 nsew signal tristate
rlabel metal2 s 389426 -960 389538 480 8 la_data_out[74]
port 370 nsew signal tristate
rlabel metal2 s 393014 -960 393126 480 8 la_data_out[75]
port 371 nsew signal tristate
rlabel metal2 s 396510 -960 396622 480 8 la_data_out[76]
port 372 nsew signal tristate
rlabel metal2 s 400098 -960 400210 480 8 la_data_out[77]
port 373 nsew signal tristate
rlabel metal2 s 403594 -960 403706 480 8 la_data_out[78]
port 374 nsew signal tristate
rlabel metal2 s 407182 -960 407294 480 8 la_data_out[79]
port 375 nsew signal tristate
rlabel metal2 s 151790 -960 151902 480 8 la_data_out[7]
port 376 nsew signal tristate
rlabel metal2 s 410770 -960 410882 480 8 la_data_out[80]
port 377 nsew signal tristate
rlabel metal2 s 414266 -960 414378 480 8 la_data_out[81]
port 378 nsew signal tristate
rlabel metal2 s 417854 -960 417966 480 8 la_data_out[82]
port 379 nsew signal tristate
rlabel metal2 s 421350 -960 421462 480 8 la_data_out[83]
port 380 nsew signal tristate
rlabel metal2 s 424938 -960 425050 480 8 la_data_out[84]
port 381 nsew signal tristate
rlabel metal2 s 428434 -960 428546 480 8 la_data_out[85]
port 382 nsew signal tristate
rlabel metal2 s 432022 -960 432134 480 8 la_data_out[86]
port 383 nsew signal tristate
rlabel metal2 s 435518 -960 435630 480 8 la_data_out[87]
port 384 nsew signal tristate
rlabel metal2 s 439106 -960 439218 480 8 la_data_out[88]
port 385 nsew signal tristate
rlabel metal2 s 442602 -960 442714 480 8 la_data_out[89]
port 386 nsew signal tristate
rlabel metal2 s 155378 -960 155490 480 8 la_data_out[8]
port 387 nsew signal tristate
rlabel metal2 s 446190 -960 446302 480 8 la_data_out[90]
port 388 nsew signal tristate
rlabel metal2 s 449778 -960 449890 480 8 la_data_out[91]
port 389 nsew signal tristate
rlabel metal2 s 453274 -960 453386 480 8 la_data_out[92]
port 390 nsew signal tristate
rlabel metal2 s 456862 -960 456974 480 8 la_data_out[93]
port 391 nsew signal tristate
rlabel metal2 s 460358 -960 460470 480 8 la_data_out[94]
port 392 nsew signal tristate
rlabel metal2 s 463946 -960 464058 480 8 la_data_out[95]
port 393 nsew signal tristate
rlabel metal2 s 467442 -960 467554 480 8 la_data_out[96]
port 394 nsew signal tristate
rlabel metal2 s 471030 -960 471142 480 8 la_data_out[97]
port 395 nsew signal tristate
rlabel metal2 s 474526 -960 474638 480 8 la_data_out[98]
port 396 nsew signal tristate
rlabel metal2 s 478114 -960 478226 480 8 la_data_out[99]
port 397 nsew signal tristate
rlabel metal2 s 158874 -960 158986 480 8 la_data_out[9]
port 398 nsew signal tristate
rlabel metal2 s 128146 -960 128258 480 8 la_oenb[0]
port 399 nsew signal input
rlabel metal2 s 482806 -960 482918 480 8 la_oenb[100]
port 400 nsew signal input
rlabel metal2 s 486394 -960 486506 480 8 la_oenb[101]
port 401 nsew signal input
rlabel metal2 s 489890 -960 490002 480 8 la_oenb[102]
port 402 nsew signal input
rlabel metal2 s 493478 -960 493590 480 8 la_oenb[103]
port 403 nsew signal input
rlabel metal2 s 497066 -960 497178 480 8 la_oenb[104]
port 404 nsew signal input
rlabel metal2 s 500562 -960 500674 480 8 la_oenb[105]
port 405 nsew signal input
rlabel metal2 s 504150 -960 504262 480 8 la_oenb[106]
port 406 nsew signal input
rlabel metal2 s 507646 -960 507758 480 8 la_oenb[107]
port 407 nsew signal input
rlabel metal2 s 511234 -960 511346 480 8 la_oenb[108]
port 408 nsew signal input
rlabel metal2 s 514730 -960 514842 480 8 la_oenb[109]
port 409 nsew signal input
rlabel metal2 s 163658 -960 163770 480 8 la_oenb[10]
port 410 nsew signal input
rlabel metal2 s 518318 -960 518430 480 8 la_oenb[110]
port 411 nsew signal input
rlabel metal2 s 521814 -960 521926 480 8 la_oenb[111]
port 412 nsew signal input
rlabel metal2 s 525402 -960 525514 480 8 la_oenb[112]
port 413 nsew signal input
rlabel metal2 s 528990 -960 529102 480 8 la_oenb[113]
port 414 nsew signal input
rlabel metal2 s 532486 -960 532598 480 8 la_oenb[114]
port 415 nsew signal input
rlabel metal2 s 536074 -960 536186 480 8 la_oenb[115]
port 416 nsew signal input
rlabel metal2 s 539570 -960 539682 480 8 la_oenb[116]
port 417 nsew signal input
rlabel metal2 s 543158 -960 543270 480 8 la_oenb[117]
port 418 nsew signal input
rlabel metal2 s 546654 -960 546766 480 8 la_oenb[118]
port 419 nsew signal input
rlabel metal2 s 550242 -960 550354 480 8 la_oenb[119]
port 420 nsew signal input
rlabel metal2 s 167154 -960 167266 480 8 la_oenb[11]
port 421 nsew signal input
rlabel metal2 s 553738 -960 553850 480 8 la_oenb[120]
port 422 nsew signal input
rlabel metal2 s 557326 -960 557438 480 8 la_oenb[121]
port 423 nsew signal input
rlabel metal2 s 560822 -960 560934 480 8 la_oenb[122]
port 424 nsew signal input
rlabel metal2 s 564410 -960 564522 480 8 la_oenb[123]
port 425 nsew signal input
rlabel metal2 s 567998 -960 568110 480 8 la_oenb[124]
port 426 nsew signal input
rlabel metal2 s 571494 -960 571606 480 8 la_oenb[125]
port 427 nsew signal input
rlabel metal2 s 575082 -960 575194 480 8 la_oenb[126]
port 428 nsew signal input
rlabel metal2 s 578578 -960 578690 480 8 la_oenb[127]
port 429 nsew signal input
rlabel metal2 s 170742 -960 170854 480 8 la_oenb[12]
port 430 nsew signal input
rlabel metal2 s 174238 -960 174350 480 8 la_oenb[13]
port 431 nsew signal input
rlabel metal2 s 177826 -960 177938 480 8 la_oenb[14]
port 432 nsew signal input
rlabel metal2 s 181414 -960 181526 480 8 la_oenb[15]
port 433 nsew signal input
rlabel metal2 s 184910 -960 185022 480 8 la_oenb[16]
port 434 nsew signal input
rlabel metal2 s 188498 -960 188610 480 8 la_oenb[17]
port 435 nsew signal input
rlabel metal2 s 191994 -960 192106 480 8 la_oenb[18]
port 436 nsew signal input
rlabel metal2 s 195582 -960 195694 480 8 la_oenb[19]
port 437 nsew signal input
rlabel metal2 s 131734 -960 131846 480 8 la_oenb[1]
port 438 nsew signal input
rlabel metal2 s 199078 -960 199190 480 8 la_oenb[20]
port 439 nsew signal input
rlabel metal2 s 202666 -960 202778 480 8 la_oenb[21]
port 440 nsew signal input
rlabel metal2 s 206162 -960 206274 480 8 la_oenb[22]
port 441 nsew signal input
rlabel metal2 s 209750 -960 209862 480 8 la_oenb[23]
port 442 nsew signal input
rlabel metal2 s 213338 -960 213450 480 8 la_oenb[24]
port 443 nsew signal input
rlabel metal2 s 216834 -960 216946 480 8 la_oenb[25]
port 444 nsew signal input
rlabel metal2 s 220422 -960 220534 480 8 la_oenb[26]
port 445 nsew signal input
rlabel metal2 s 223918 -960 224030 480 8 la_oenb[27]
port 446 nsew signal input
rlabel metal2 s 227506 -960 227618 480 8 la_oenb[28]
port 447 nsew signal input
rlabel metal2 s 231002 -960 231114 480 8 la_oenb[29]
port 448 nsew signal input
rlabel metal2 s 135230 -960 135342 480 8 la_oenb[2]
port 449 nsew signal input
rlabel metal2 s 234590 -960 234702 480 8 la_oenb[30]
port 450 nsew signal input
rlabel metal2 s 238086 -960 238198 480 8 la_oenb[31]
port 451 nsew signal input
rlabel metal2 s 241674 -960 241786 480 8 la_oenb[32]
port 452 nsew signal input
rlabel metal2 s 245170 -960 245282 480 8 la_oenb[33]
port 453 nsew signal input
rlabel metal2 s 248758 -960 248870 480 8 la_oenb[34]
port 454 nsew signal input
rlabel metal2 s 252346 -960 252458 480 8 la_oenb[35]
port 455 nsew signal input
rlabel metal2 s 255842 -960 255954 480 8 la_oenb[36]
port 456 nsew signal input
rlabel metal2 s 259430 -960 259542 480 8 la_oenb[37]
port 457 nsew signal input
rlabel metal2 s 262926 -960 263038 480 8 la_oenb[38]
port 458 nsew signal input
rlabel metal2 s 266514 -960 266626 480 8 la_oenb[39]
port 459 nsew signal input
rlabel metal2 s 138818 -960 138930 480 8 la_oenb[3]
port 460 nsew signal input
rlabel metal2 s 270010 -960 270122 480 8 la_oenb[40]
port 461 nsew signal input
rlabel metal2 s 273598 -960 273710 480 8 la_oenb[41]
port 462 nsew signal input
rlabel metal2 s 277094 -960 277206 480 8 la_oenb[42]
port 463 nsew signal input
rlabel metal2 s 280682 -960 280794 480 8 la_oenb[43]
port 464 nsew signal input
rlabel metal2 s 284270 -960 284382 480 8 la_oenb[44]
port 465 nsew signal input
rlabel metal2 s 287766 -960 287878 480 8 la_oenb[45]
port 466 nsew signal input
rlabel metal2 s 291354 -960 291466 480 8 la_oenb[46]
port 467 nsew signal input
rlabel metal2 s 294850 -960 294962 480 8 la_oenb[47]
port 468 nsew signal input
rlabel metal2 s 298438 -960 298550 480 8 la_oenb[48]
port 469 nsew signal input
rlabel metal2 s 301934 -960 302046 480 8 la_oenb[49]
port 470 nsew signal input
rlabel metal2 s 142406 -960 142518 480 8 la_oenb[4]
port 471 nsew signal input
rlabel metal2 s 305522 -960 305634 480 8 la_oenb[50]
port 472 nsew signal input
rlabel metal2 s 309018 -960 309130 480 8 la_oenb[51]
port 473 nsew signal input
rlabel metal2 s 312606 -960 312718 480 8 la_oenb[52]
port 474 nsew signal input
rlabel metal2 s 316194 -960 316306 480 8 la_oenb[53]
port 475 nsew signal input
rlabel metal2 s 319690 -960 319802 480 8 la_oenb[54]
port 476 nsew signal input
rlabel metal2 s 323278 -960 323390 480 8 la_oenb[55]
port 477 nsew signal input
rlabel metal2 s 326774 -960 326886 480 8 la_oenb[56]
port 478 nsew signal input
rlabel metal2 s 330362 -960 330474 480 8 la_oenb[57]
port 479 nsew signal input
rlabel metal2 s 333858 -960 333970 480 8 la_oenb[58]
port 480 nsew signal input
rlabel metal2 s 337446 -960 337558 480 8 la_oenb[59]
port 481 nsew signal input
rlabel metal2 s 145902 -960 146014 480 8 la_oenb[5]
port 482 nsew signal input
rlabel metal2 s 340942 -960 341054 480 8 la_oenb[60]
port 483 nsew signal input
rlabel metal2 s 344530 -960 344642 480 8 la_oenb[61]
port 484 nsew signal input
rlabel metal2 s 348026 -960 348138 480 8 la_oenb[62]
port 485 nsew signal input
rlabel metal2 s 351614 -960 351726 480 8 la_oenb[63]
port 486 nsew signal input
rlabel metal2 s 355202 -960 355314 480 8 la_oenb[64]
port 487 nsew signal input
rlabel metal2 s 358698 -960 358810 480 8 la_oenb[65]
port 488 nsew signal input
rlabel metal2 s 362286 -960 362398 480 8 la_oenb[66]
port 489 nsew signal input
rlabel metal2 s 365782 -960 365894 480 8 la_oenb[67]
port 490 nsew signal input
rlabel metal2 s 369370 -960 369482 480 8 la_oenb[68]
port 491 nsew signal input
rlabel metal2 s 372866 -960 372978 480 8 la_oenb[69]
port 492 nsew signal input
rlabel metal2 s 149490 -960 149602 480 8 la_oenb[6]
port 493 nsew signal input
rlabel metal2 s 376454 -960 376566 480 8 la_oenb[70]
port 494 nsew signal input
rlabel metal2 s 379950 -960 380062 480 8 la_oenb[71]
port 495 nsew signal input
rlabel metal2 s 383538 -960 383650 480 8 la_oenb[72]
port 496 nsew signal input
rlabel metal2 s 387126 -960 387238 480 8 la_oenb[73]
port 497 nsew signal input
rlabel metal2 s 390622 -960 390734 480 8 la_oenb[74]
port 498 nsew signal input
rlabel metal2 s 394210 -960 394322 480 8 la_oenb[75]
port 499 nsew signal input
rlabel metal2 s 397706 -960 397818 480 8 la_oenb[76]
port 500 nsew signal input
rlabel metal2 s 401294 -960 401406 480 8 la_oenb[77]
port 501 nsew signal input
rlabel metal2 s 404790 -960 404902 480 8 la_oenb[78]
port 502 nsew signal input
rlabel metal2 s 408378 -960 408490 480 8 la_oenb[79]
port 503 nsew signal input
rlabel metal2 s 152986 -960 153098 480 8 la_oenb[7]
port 504 nsew signal input
rlabel metal2 s 411874 -960 411986 480 8 la_oenb[80]
port 505 nsew signal input
rlabel metal2 s 415462 -960 415574 480 8 la_oenb[81]
port 506 nsew signal input
rlabel metal2 s 418958 -960 419070 480 8 la_oenb[82]
port 507 nsew signal input
rlabel metal2 s 422546 -960 422658 480 8 la_oenb[83]
port 508 nsew signal input
rlabel metal2 s 426134 -960 426246 480 8 la_oenb[84]
port 509 nsew signal input
rlabel metal2 s 429630 -960 429742 480 8 la_oenb[85]
port 510 nsew signal input
rlabel metal2 s 433218 -960 433330 480 8 la_oenb[86]
port 511 nsew signal input
rlabel metal2 s 436714 -960 436826 480 8 la_oenb[87]
port 512 nsew signal input
rlabel metal2 s 440302 -960 440414 480 8 la_oenb[88]
port 513 nsew signal input
rlabel metal2 s 443798 -960 443910 480 8 la_oenb[89]
port 514 nsew signal input
rlabel metal2 s 156574 -960 156686 480 8 la_oenb[8]
port 515 nsew signal input
rlabel metal2 s 447386 -960 447498 480 8 la_oenb[90]
port 516 nsew signal input
rlabel metal2 s 450882 -960 450994 480 8 la_oenb[91]
port 517 nsew signal input
rlabel metal2 s 454470 -960 454582 480 8 la_oenb[92]
port 518 nsew signal input
rlabel metal2 s 458058 -960 458170 480 8 la_oenb[93]
port 519 nsew signal input
rlabel metal2 s 461554 -960 461666 480 8 la_oenb[94]
port 520 nsew signal input
rlabel metal2 s 465142 -960 465254 480 8 la_oenb[95]
port 521 nsew signal input
rlabel metal2 s 468638 -960 468750 480 8 la_oenb[96]
port 522 nsew signal input
rlabel metal2 s 472226 -960 472338 480 8 la_oenb[97]
port 523 nsew signal input
rlabel metal2 s 475722 -960 475834 480 8 la_oenb[98]
port 524 nsew signal input
rlabel metal2 s 479310 -960 479422 480 8 la_oenb[99]
port 525 nsew signal input
rlabel metal2 s 160070 -960 160182 480 8 la_oenb[9]
port 526 nsew signal input
rlabel metal2 s 579774 -960 579886 480 8 user_clock2
port 527 nsew signal input
rlabel metal2 s 580970 -960 581082 480 8 user_irq[0]
port 528 nsew signal tristate
rlabel metal2 s 582166 -960 582278 480 8 user_irq[1]
port 529 nsew signal tristate
rlabel metal2 s 583362 -960 583474 480 8 user_irq[2]
port 530 nsew signal tristate
rlabel metal5 s -2006 -934 585930 -314 8 vccd1
port 531 nsew power input
rlabel metal5 s -2966 1876 586890 2476 6 vccd1
port 531 nsew power input
rlabel metal5 s -2966 37876 586890 38476 6 vccd1
port 531 nsew power input
rlabel metal5 s -2966 73876 586890 74476 6 vccd1
port 531 nsew power input
rlabel metal5 s -2966 109876 586890 110476 6 vccd1
port 531 nsew power input
rlabel metal5 s -2966 145876 586890 146476 6 vccd1
port 531 nsew power input
rlabel metal5 s -2966 181876 586890 182476 6 vccd1
port 531 nsew power input
rlabel metal5 s -2966 217876 586890 218476 6 vccd1
port 531 nsew power input
rlabel metal5 s -2966 253876 586890 254476 6 vccd1
port 531 nsew power input
rlabel metal5 s -2966 289876 586890 290476 6 vccd1
port 531 nsew power input
rlabel metal5 s -2966 325876 586890 326476 6 vccd1
port 531 nsew power input
rlabel metal5 s -2966 361876 586890 362476 6 vccd1
port 531 nsew power input
rlabel metal5 s -2966 397876 586890 398476 6 vccd1
port 531 nsew power input
rlabel metal5 s -2966 433876 586890 434476 6 vccd1
port 531 nsew power input
rlabel metal5 s -2966 469876 586890 470476 6 vccd1
port 531 nsew power input
rlabel metal5 s -2966 505876 586890 506476 6 vccd1
port 531 nsew power input
rlabel metal5 s -2966 541876 586890 542476 6 vccd1
port 531 nsew power input
rlabel metal5 s -2966 577876 586890 578476 6 vccd1
port 531 nsew power input
rlabel metal5 s -2966 613876 586890 614476 6 vccd1
port 531 nsew power input
rlabel metal5 s -2966 649876 586890 650476 6 vccd1
port 531 nsew power input
rlabel metal5 s -2966 685876 586890 686476 6 vccd1
port 531 nsew power input
rlabel metal5 s -2006 704250 585930 704870 6 vccd1
port 531 nsew power input
rlabel metal4 s 72804 -1894 73404 38000 6 vccd1
port 531 nsew power input
rlabel metal4 s 108804 -1894 109404 38000 6 vccd1
port 531 nsew power input
rlabel metal4 s 144804 -1894 145404 38000 6 vccd1
port 531 nsew power input
rlabel metal4 s 180804 -1894 181404 38000 6 vccd1
port 531 nsew power input
rlabel metal4 s 216804 -1894 217404 38000 6 vccd1
port 531 nsew power input
rlabel metal4 s 72804 243568 73404 338000 6 vccd1
port 531 nsew power input
rlabel metal4 s 108804 243568 109404 338000 6 vccd1
port 531 nsew power input
rlabel metal4 s 144804 243568 145404 338000 6 vccd1
port 531 nsew power input
rlabel metal4 s 360804 -1894 361404 338000 6 vccd1
port 531 nsew power input
rlabel metal4 s 396804 -1894 397404 338000 6 vccd1
port 531 nsew power input
rlabel metal4 s 432804 -1894 433404 338000 6 vccd1
port 531 nsew power input
rlabel metal4 s 468804 -1894 469404 338000 6 vccd1
port 531 nsew power input
rlabel metal4 s -2006 -934 -1386 704870 4 vccd1
port 531 nsew power input
rlabel metal4 s 585310 -934 585930 704870 6 vccd1
port 531 nsew power input
rlabel metal4 s 804 -1894 1404 705830 6 vccd1
port 531 nsew power input
rlabel metal4 s 36804 -1894 37404 705830 6 vccd1
port 531 nsew power input
rlabel metal4 s 72804 425308 73404 705830 6 vccd1
port 531 nsew power input
rlabel metal4 s 108804 425308 109404 705830 6 vccd1
port 531 nsew power input
rlabel metal4 s 144804 425308 145404 705830 6 vccd1
port 531 nsew power input
rlabel metal4 s 180804 243568 181404 705830 6 vccd1
port 531 nsew power input
rlabel metal4 s 216804 243568 217404 705830 6 vccd1
port 531 nsew power input
rlabel metal4 s 252804 -1894 253404 705830 6 vccd1
port 531 nsew power input
rlabel metal4 s 288804 -1894 289404 705830 6 vccd1
port 531 nsew power input
rlabel metal4 s 324804 -1894 325404 705830 6 vccd1
port 531 nsew power input
rlabel metal4 s 360804 425308 361404 705830 6 vccd1
port 531 nsew power input
rlabel metal4 s 396804 425308 397404 705830 6 vccd1
port 531 nsew power input
rlabel metal4 s 432804 425308 433404 705830 6 vccd1
port 531 nsew power input
rlabel metal4 s 468804 425308 469404 705830 6 vccd1
port 531 nsew power input
rlabel metal4 s 504804 -1894 505404 705830 6 vccd1
port 531 nsew power input
rlabel metal4 s 540804 -1894 541404 705830 6 vccd1
port 531 nsew power input
rlabel metal4 s 576804 -1894 577404 705830 6 vccd1
port 531 nsew power input
rlabel metal5 s -3926 -2854 587850 -2234 8 vccd2
port 532 nsew power input
rlabel metal5 s -4886 5576 588810 6176 6 vccd2
port 532 nsew power input
rlabel metal5 s -4886 41576 588810 42176 6 vccd2
port 532 nsew power input
rlabel metal5 s -4886 77576 588810 78176 6 vccd2
port 532 nsew power input
rlabel metal5 s -4886 113576 588810 114176 6 vccd2
port 532 nsew power input
rlabel metal5 s -4886 149576 588810 150176 6 vccd2
port 532 nsew power input
rlabel metal5 s -4886 185576 588810 186176 6 vccd2
port 532 nsew power input
rlabel metal5 s -4886 221576 588810 222176 6 vccd2
port 532 nsew power input
rlabel metal5 s -4886 257576 588810 258176 6 vccd2
port 532 nsew power input
rlabel metal5 s -4886 293576 588810 294176 6 vccd2
port 532 nsew power input
rlabel metal5 s -4886 329576 588810 330176 6 vccd2
port 532 nsew power input
rlabel metal5 s -4886 365576 588810 366176 6 vccd2
port 532 nsew power input
rlabel metal5 s -4886 401576 588810 402176 6 vccd2
port 532 nsew power input
rlabel metal5 s -4886 437576 588810 438176 6 vccd2
port 532 nsew power input
rlabel metal5 s -4886 473576 588810 474176 6 vccd2
port 532 nsew power input
rlabel metal5 s -4886 509576 588810 510176 6 vccd2
port 532 nsew power input
rlabel metal5 s -4886 545576 588810 546176 6 vccd2
port 532 nsew power input
rlabel metal5 s -4886 581576 588810 582176 6 vccd2
port 532 nsew power input
rlabel metal5 s -4886 617576 588810 618176 6 vccd2
port 532 nsew power input
rlabel metal5 s -4886 653576 588810 654176 6 vccd2
port 532 nsew power input
rlabel metal5 s -4886 689576 588810 690176 6 vccd2
port 532 nsew power input
rlabel metal5 s -3926 706170 587850 706790 6 vccd2
port 532 nsew power input
rlabel metal4 s 40504 -3814 41104 38000 6 vccd2
port 532 nsew power input
rlabel metal4 s 76504 -3814 77104 38000 6 vccd2
port 532 nsew power input
rlabel metal4 s 112504 -3814 113104 38000 6 vccd2
port 532 nsew power input
rlabel metal4 s 148504 -3814 149104 38000 6 vccd2
port 532 nsew power input
rlabel metal4 s 184504 -3814 185104 38000 6 vccd2
port 532 nsew power input
rlabel metal4 s 220504 -3814 221104 38000 6 vccd2
port 532 nsew power input
rlabel metal4 s 40504 243568 41104 338000 6 vccd2
port 532 nsew power input
rlabel metal4 s 76504 243568 77104 338000 6 vccd2
port 532 nsew power input
rlabel metal4 s 112504 243568 113104 338000 6 vccd2
port 532 nsew power input
rlabel metal4 s 148504 243568 149104 338000 6 vccd2
port 532 nsew power input
rlabel metal4 s 364504 -3814 365104 338000 6 vccd2
port 532 nsew power input
rlabel metal4 s 400504 -3814 401104 338000 6 vccd2
port 532 nsew power input
rlabel metal4 s 436504 -3814 437104 338000 6 vccd2
port 532 nsew power input
rlabel metal4 s 472504 -3814 473104 338000 6 vccd2
port 532 nsew power input
rlabel metal4 s -3926 -2854 -3306 706790 4 vccd2
port 532 nsew power input
rlabel metal4 s 587230 -2854 587850 706790 6 vccd2
port 532 nsew power input
rlabel metal4 s 4504 -3814 5104 707750 6 vccd2
port 532 nsew power input
rlabel metal4 s 40504 425308 41104 707750 6 vccd2
port 532 nsew power input
rlabel metal4 s 76504 425308 77104 707750 6 vccd2
port 532 nsew power input
rlabel metal4 s 112504 425308 113104 707750 6 vccd2
port 532 nsew power input
rlabel metal4 s 148504 425308 149104 707750 6 vccd2
port 532 nsew power input
rlabel metal4 s 184504 243568 185104 707750 6 vccd2
port 532 nsew power input
rlabel metal4 s 220504 243568 221104 707750 6 vccd2
port 532 nsew power input
rlabel metal4 s 256504 -3814 257104 707750 6 vccd2
port 532 nsew power input
rlabel metal4 s 292504 -3814 293104 707750 6 vccd2
port 532 nsew power input
rlabel metal4 s 328504 -3814 329104 707750 6 vccd2
port 532 nsew power input
rlabel metal4 s 364504 425308 365104 707750 6 vccd2
port 532 nsew power input
rlabel metal4 s 400504 425308 401104 707750 6 vccd2
port 532 nsew power input
rlabel metal4 s 436504 425308 437104 707750 6 vccd2
port 532 nsew power input
rlabel metal4 s 472504 425308 473104 707750 6 vccd2
port 532 nsew power input
rlabel metal4 s 508504 -3814 509104 707750 6 vccd2
port 532 nsew power input
rlabel metal4 s 544504 -3814 545104 707750 6 vccd2
port 532 nsew power input
rlabel metal4 s 580504 -3814 581104 707750 6 vccd2
port 532 nsew power input
rlabel metal5 s -5846 -4774 589770 -4154 8 vdda1
port 533 nsew power input
rlabel metal5 s -6806 9276 590730 9876 6 vdda1
port 533 nsew power input
rlabel metal5 s -6806 45276 590730 45876 6 vdda1
port 533 nsew power input
rlabel metal5 s -6806 81276 590730 81876 6 vdda1
port 533 nsew power input
rlabel metal5 s -6806 117276 590730 117876 6 vdda1
port 533 nsew power input
rlabel metal5 s -6806 153276 590730 153876 6 vdda1
port 533 nsew power input
rlabel metal5 s -6806 189276 590730 189876 6 vdda1
port 533 nsew power input
rlabel metal5 s -6806 225276 590730 225876 6 vdda1
port 533 nsew power input
rlabel metal5 s -6806 261276 590730 261876 6 vdda1
port 533 nsew power input
rlabel metal5 s -6806 297276 590730 297876 6 vdda1
port 533 nsew power input
rlabel metal5 s -6806 333276 590730 333876 6 vdda1
port 533 nsew power input
rlabel metal5 s -6806 369276 590730 369876 6 vdda1
port 533 nsew power input
rlabel metal5 s -6806 405276 590730 405876 6 vdda1
port 533 nsew power input
rlabel metal5 s -6806 441276 590730 441876 6 vdda1
port 533 nsew power input
rlabel metal5 s -6806 477276 590730 477876 6 vdda1
port 533 nsew power input
rlabel metal5 s -6806 513276 590730 513876 6 vdda1
port 533 nsew power input
rlabel metal5 s -6806 549276 590730 549876 6 vdda1
port 533 nsew power input
rlabel metal5 s -6806 585276 590730 585876 6 vdda1
port 533 nsew power input
rlabel metal5 s -6806 621276 590730 621876 6 vdda1
port 533 nsew power input
rlabel metal5 s -6806 657276 590730 657876 6 vdda1
port 533 nsew power input
rlabel metal5 s -6806 693276 590730 693876 6 vdda1
port 533 nsew power input
rlabel metal5 s -5846 708090 589770 708710 6 vdda1
port 533 nsew power input
rlabel metal4 s 44204 -5734 44804 38000 6 vdda1
port 533 nsew power input
rlabel metal4 s 80204 -5734 80804 38000 6 vdda1
port 533 nsew power input
rlabel metal4 s 116204 -5734 116804 38000 6 vdda1
port 533 nsew power input
rlabel metal4 s 152204 -5734 152804 38000 6 vdda1
port 533 nsew power input
rlabel metal4 s 188204 -5734 188804 38000 6 vdda1
port 533 nsew power input
rlabel metal4 s 224204 -5734 224804 38000 6 vdda1
port 533 nsew power input
rlabel metal4 s 44204 243568 44804 338000 6 vdda1
port 533 nsew power input
rlabel metal4 s 80204 243568 80804 338000 6 vdda1
port 533 nsew power input
rlabel metal4 s 116204 243568 116804 338000 6 vdda1
port 533 nsew power input
rlabel metal4 s 152204 243568 152804 338000 6 vdda1
port 533 nsew power input
rlabel metal4 s 368204 -5734 368804 338000 6 vdda1
port 533 nsew power input
rlabel metal4 s 404204 -5734 404804 338000 6 vdda1
port 533 nsew power input
rlabel metal4 s 440204 -5734 440804 338000 6 vdda1
port 533 nsew power input
rlabel metal4 s 476204 -5734 476804 338000 6 vdda1
port 533 nsew power input
rlabel metal4 s -5846 -4774 -5226 708710 4 vdda1
port 533 nsew power input
rlabel metal4 s 589150 -4774 589770 708710 6 vdda1
port 533 nsew power input
rlabel metal4 s 8204 -5734 8804 709670 6 vdda1
port 533 nsew power input
rlabel metal4 s 44204 425308 44804 709670 6 vdda1
port 533 nsew power input
rlabel metal4 s 80204 425308 80804 709670 6 vdda1
port 533 nsew power input
rlabel metal4 s 116204 425308 116804 709670 6 vdda1
port 533 nsew power input
rlabel metal4 s 152204 425308 152804 709670 6 vdda1
port 533 nsew power input
rlabel metal4 s 188204 243568 188804 709670 6 vdda1
port 533 nsew power input
rlabel metal4 s 224204 243568 224804 709670 6 vdda1
port 533 nsew power input
rlabel metal4 s 260204 -5734 260804 709670 6 vdda1
port 533 nsew power input
rlabel metal4 s 296204 -5734 296804 709670 6 vdda1
port 533 nsew power input
rlabel metal4 s 332204 -5734 332804 709670 6 vdda1
port 533 nsew power input
rlabel metal4 s 368204 425308 368804 709670 6 vdda1
port 533 nsew power input
rlabel metal4 s 404204 425308 404804 709670 6 vdda1
port 533 nsew power input
rlabel metal4 s 440204 425308 440804 709670 6 vdda1
port 533 nsew power input
rlabel metal4 s 476204 425308 476804 709670 6 vdda1
port 533 nsew power input
rlabel metal4 s 512204 -5734 512804 709670 6 vdda1
port 533 nsew power input
rlabel metal4 s 548204 -5734 548804 709670 6 vdda1
port 533 nsew power input
rlabel metal5 s -7766 -6694 591690 -6074 8 vdda2
port 534 nsew power input
rlabel metal5 s -8726 12976 592650 13576 6 vdda2
port 534 nsew power input
rlabel metal5 s -8726 48976 592650 49576 6 vdda2
port 534 nsew power input
rlabel metal5 s -8726 84976 592650 85576 6 vdda2
port 534 nsew power input
rlabel metal5 s -8726 120976 592650 121576 6 vdda2
port 534 nsew power input
rlabel metal5 s -8726 156976 592650 157576 6 vdda2
port 534 nsew power input
rlabel metal5 s -8726 192976 592650 193576 6 vdda2
port 534 nsew power input
rlabel metal5 s -8726 228976 592650 229576 6 vdda2
port 534 nsew power input
rlabel metal5 s -8726 264976 592650 265576 6 vdda2
port 534 nsew power input
rlabel metal5 s -8726 300976 592650 301576 6 vdda2
port 534 nsew power input
rlabel metal5 s -8726 336976 592650 337576 6 vdda2
port 534 nsew power input
rlabel metal5 s -8726 372976 592650 373576 6 vdda2
port 534 nsew power input
rlabel metal5 s -8726 408976 592650 409576 6 vdda2
port 534 nsew power input
rlabel metal5 s -8726 444976 592650 445576 6 vdda2
port 534 nsew power input
rlabel metal5 s -8726 480976 592650 481576 6 vdda2
port 534 nsew power input
rlabel metal5 s -8726 516976 592650 517576 6 vdda2
port 534 nsew power input
rlabel metal5 s -8726 552976 592650 553576 6 vdda2
port 534 nsew power input
rlabel metal5 s -8726 588976 592650 589576 6 vdda2
port 534 nsew power input
rlabel metal5 s -8726 624976 592650 625576 6 vdda2
port 534 nsew power input
rlabel metal5 s -8726 660976 592650 661576 6 vdda2
port 534 nsew power input
rlabel metal5 s -8726 696976 592650 697576 6 vdda2
port 534 nsew power input
rlabel metal5 s -7766 710010 591690 710630 6 vdda2
port 534 nsew power input
rlabel metal4 s 47904 -7654 48504 38000 6 vdda2
port 534 nsew power input
rlabel metal4 s 83904 -7654 84504 38000 6 vdda2
port 534 nsew power input
rlabel metal4 s 119904 -7654 120504 38000 6 vdda2
port 534 nsew power input
rlabel metal4 s 155904 -7654 156504 38000 6 vdda2
port 534 nsew power input
rlabel metal4 s 191904 -7654 192504 38000 6 vdda2
port 534 nsew power input
rlabel metal4 s 227904 -7654 228504 38000 6 vdda2
port 534 nsew power input
rlabel metal4 s 47904 243568 48504 338000 6 vdda2
port 534 nsew power input
rlabel metal4 s 83904 243568 84504 338000 6 vdda2
port 534 nsew power input
rlabel metal4 s 119904 243568 120504 338000 6 vdda2
port 534 nsew power input
rlabel metal4 s 155904 243568 156504 338000 6 vdda2
port 534 nsew power input
rlabel metal4 s 371904 -7654 372504 338000 6 vdda2
port 534 nsew power input
rlabel metal4 s 407904 -7654 408504 338000 6 vdda2
port 534 nsew power input
rlabel metal4 s 443904 -7654 444504 338000 6 vdda2
port 534 nsew power input
rlabel metal4 s -7766 -6694 -7146 710630 4 vdda2
port 534 nsew power input
rlabel metal4 s 591070 -6694 591690 710630 6 vdda2
port 534 nsew power input
rlabel metal4 s 11904 -7654 12504 711590 6 vdda2
port 534 nsew power input
rlabel metal4 s 47904 425308 48504 711590 6 vdda2
port 534 nsew power input
rlabel metal4 s 83904 425308 84504 711590 6 vdda2
port 534 nsew power input
rlabel metal4 s 119904 425308 120504 711590 6 vdda2
port 534 nsew power input
rlabel metal4 s 155904 425308 156504 711590 6 vdda2
port 534 nsew power input
rlabel metal4 s 191904 243568 192504 711590 6 vdda2
port 534 nsew power input
rlabel metal4 s 227904 243568 228504 711590 6 vdda2
port 534 nsew power input
rlabel metal4 s 263904 -7654 264504 711590 6 vdda2
port 534 nsew power input
rlabel metal4 s 299904 -7654 300504 711590 6 vdda2
port 534 nsew power input
rlabel metal4 s 335904 -7654 336504 711590 6 vdda2
port 534 nsew power input
rlabel metal4 s 371904 425308 372504 711590 6 vdda2
port 534 nsew power input
rlabel metal4 s 407904 425308 408504 711590 6 vdda2
port 534 nsew power input
rlabel metal4 s 443904 425308 444504 711590 6 vdda2
port 534 nsew power input
rlabel metal4 s 479904 -7654 480504 711590 6 vdda2
port 534 nsew power input
rlabel metal4 s 515904 -7654 516504 711590 6 vdda2
port 534 nsew power input
rlabel metal4 s 551904 -7654 552504 711590 6 vdda2
port 534 nsew power input
rlabel metal5 s -6806 -5734 590730 -5114 8 vssa1
port 535 nsew ground input
rlabel metal5 s -6806 27276 590730 27876 6 vssa1
port 535 nsew ground input
rlabel metal5 s -6806 63276 590730 63876 6 vssa1
port 535 nsew ground input
rlabel metal5 s -6806 99276 590730 99876 6 vssa1
port 535 nsew ground input
rlabel metal5 s -6806 135276 590730 135876 6 vssa1
port 535 nsew ground input
rlabel metal5 s -6806 171276 590730 171876 6 vssa1
port 535 nsew ground input
rlabel metal5 s -6806 207276 590730 207876 6 vssa1
port 535 nsew ground input
rlabel metal5 s -6806 243276 590730 243876 6 vssa1
port 535 nsew ground input
rlabel metal5 s -6806 279276 590730 279876 6 vssa1
port 535 nsew ground input
rlabel metal5 s -6806 315276 590730 315876 6 vssa1
port 535 nsew ground input
rlabel metal5 s -6806 351276 590730 351876 6 vssa1
port 535 nsew ground input
rlabel metal5 s -6806 387276 590730 387876 6 vssa1
port 535 nsew ground input
rlabel metal5 s -6806 423276 590730 423876 6 vssa1
port 535 nsew ground input
rlabel metal5 s -6806 459276 590730 459876 6 vssa1
port 535 nsew ground input
rlabel metal5 s -6806 495276 590730 495876 6 vssa1
port 535 nsew ground input
rlabel metal5 s -6806 531276 590730 531876 6 vssa1
port 535 nsew ground input
rlabel metal5 s -6806 567276 590730 567876 6 vssa1
port 535 nsew ground input
rlabel metal5 s -6806 603276 590730 603876 6 vssa1
port 535 nsew ground input
rlabel metal5 s -6806 639276 590730 639876 6 vssa1
port 535 nsew ground input
rlabel metal5 s -6806 675276 590730 675876 6 vssa1
port 535 nsew ground input
rlabel metal5 s -6806 709050 590730 709670 6 vssa1
port 535 nsew ground input
rlabel metal4 s 62204 -5734 62804 38000 6 vssa1
port 535 nsew ground input
rlabel metal4 s 98204 -5734 98804 38000 6 vssa1
port 535 nsew ground input
rlabel metal4 s 134204 -5734 134804 38000 6 vssa1
port 535 nsew ground input
rlabel metal4 s 170204 -5734 170804 38000 6 vssa1
port 535 nsew ground input
rlabel metal4 s 206204 -5734 206804 38000 6 vssa1
port 535 nsew ground input
rlabel metal4 s 62204 243568 62804 338000 6 vssa1
port 535 nsew ground input
rlabel metal4 s 98204 243568 98804 338000 6 vssa1
port 535 nsew ground input
rlabel metal4 s 134204 243568 134804 338000 6 vssa1
port 535 nsew ground input
rlabel metal4 s 170204 243568 170804 338000 6 vssa1
port 535 nsew ground input
rlabel metal4 s 350204 -5734 350804 338000 6 vssa1
port 535 nsew ground input
rlabel metal4 s 386204 -5734 386804 338000 6 vssa1
port 535 nsew ground input
rlabel metal4 s 422204 -5734 422804 338000 6 vssa1
port 535 nsew ground input
rlabel metal4 s 458204 -5734 458804 338000 6 vssa1
port 535 nsew ground input
rlabel metal4 s -6806 -5734 -6186 709670 4 vssa1
port 535 nsew ground input
rlabel metal4 s 26204 -5734 26804 709670 6 vssa1
port 535 nsew ground input
rlabel metal4 s 62204 425308 62804 709670 6 vssa1
port 535 nsew ground input
rlabel metal4 s 98204 425308 98804 709670 6 vssa1
port 535 nsew ground input
rlabel metal4 s 134204 425308 134804 709670 6 vssa1
port 535 nsew ground input
rlabel metal4 s 170204 425308 170804 709670 6 vssa1
port 535 nsew ground input
rlabel metal4 s 206204 243568 206804 709670 6 vssa1
port 535 nsew ground input
rlabel metal4 s 242204 -5734 242804 709670 6 vssa1
port 535 nsew ground input
rlabel metal4 s 278204 -5734 278804 709670 6 vssa1
port 535 nsew ground input
rlabel metal4 s 314204 -5734 314804 709670 6 vssa1
port 535 nsew ground input
rlabel metal4 s 350204 425308 350804 709670 6 vssa1
port 535 nsew ground input
rlabel metal4 s 386204 425308 386804 709670 6 vssa1
port 535 nsew ground input
rlabel metal4 s 422204 425308 422804 709670 6 vssa1
port 535 nsew ground input
rlabel metal4 s 458204 425308 458804 709670 6 vssa1
port 535 nsew ground input
rlabel metal4 s 494204 -5734 494804 709670 6 vssa1
port 535 nsew ground input
rlabel metal4 s 530204 -5734 530804 709670 6 vssa1
port 535 nsew ground input
rlabel metal4 s 566204 -5734 566804 709670 6 vssa1
port 535 nsew ground input
rlabel metal4 s 590110 -5734 590730 709670 6 vssa1
port 535 nsew ground input
rlabel metal5 s -8726 -7654 592650 -7034 8 vssa2
port 536 nsew ground input
rlabel metal5 s -8726 30976 592650 31576 6 vssa2
port 536 nsew ground input
rlabel metal5 s -8726 66976 592650 67576 6 vssa2
port 536 nsew ground input
rlabel metal5 s -8726 102976 592650 103576 6 vssa2
port 536 nsew ground input
rlabel metal5 s -8726 138976 592650 139576 6 vssa2
port 536 nsew ground input
rlabel metal5 s -8726 174976 592650 175576 6 vssa2
port 536 nsew ground input
rlabel metal5 s -8726 210976 592650 211576 6 vssa2
port 536 nsew ground input
rlabel metal5 s -8726 246976 592650 247576 6 vssa2
port 536 nsew ground input
rlabel metal5 s -8726 282976 592650 283576 6 vssa2
port 536 nsew ground input
rlabel metal5 s -8726 318976 592650 319576 6 vssa2
port 536 nsew ground input
rlabel metal5 s -8726 354976 592650 355576 6 vssa2
port 536 nsew ground input
rlabel metal5 s -8726 390976 592650 391576 6 vssa2
port 536 nsew ground input
rlabel metal5 s -8726 426976 592650 427576 6 vssa2
port 536 nsew ground input
rlabel metal5 s -8726 462976 592650 463576 6 vssa2
port 536 nsew ground input
rlabel metal5 s -8726 498976 592650 499576 6 vssa2
port 536 nsew ground input
rlabel metal5 s -8726 534976 592650 535576 6 vssa2
port 536 nsew ground input
rlabel metal5 s -8726 570976 592650 571576 6 vssa2
port 536 nsew ground input
rlabel metal5 s -8726 606976 592650 607576 6 vssa2
port 536 nsew ground input
rlabel metal5 s -8726 642976 592650 643576 6 vssa2
port 536 nsew ground input
rlabel metal5 s -8726 678976 592650 679576 6 vssa2
port 536 nsew ground input
rlabel metal5 s -8726 710970 592650 711590 6 vssa2
port 536 nsew ground input
rlabel metal4 s 65904 -7654 66504 38000 6 vssa2
port 536 nsew ground input
rlabel metal4 s 101904 -7654 102504 38000 6 vssa2
port 536 nsew ground input
rlabel metal4 s 137904 -7654 138504 38000 6 vssa2
port 536 nsew ground input
rlabel metal4 s 173904 -7654 174504 38000 6 vssa2
port 536 nsew ground input
rlabel metal4 s 209904 -7654 210504 38000 6 vssa2
port 536 nsew ground input
rlabel metal4 s 65904 243568 66504 338000 6 vssa2
port 536 nsew ground input
rlabel metal4 s 101904 243568 102504 338000 6 vssa2
port 536 nsew ground input
rlabel metal4 s 137904 243568 138504 338000 6 vssa2
port 536 nsew ground input
rlabel metal4 s 173904 243568 174504 338000 6 vssa2
port 536 nsew ground input
rlabel metal4 s 353904 -7654 354504 338000 6 vssa2
port 536 nsew ground input
rlabel metal4 s 389904 -7654 390504 338000 6 vssa2
port 536 nsew ground input
rlabel metal4 s 425904 -7654 426504 338000 6 vssa2
port 536 nsew ground input
rlabel metal4 s 461904 -7654 462504 338000 6 vssa2
port 536 nsew ground input
rlabel metal4 s -8726 -7654 -8106 711590 4 vssa2
port 536 nsew ground input
rlabel metal4 s 29904 -7654 30504 711590 6 vssa2
port 536 nsew ground input
rlabel metal4 s 65904 425308 66504 711590 6 vssa2
port 536 nsew ground input
rlabel metal4 s 101904 425308 102504 711590 6 vssa2
port 536 nsew ground input
rlabel metal4 s 137904 425308 138504 711590 6 vssa2
port 536 nsew ground input
rlabel metal4 s 173904 425308 174504 711590 6 vssa2
port 536 nsew ground input
rlabel metal4 s 209904 243568 210504 711590 6 vssa2
port 536 nsew ground input
rlabel metal4 s 245904 -7654 246504 711590 6 vssa2
port 536 nsew ground input
rlabel metal4 s 281904 -7654 282504 711590 6 vssa2
port 536 nsew ground input
rlabel metal4 s 317904 -7654 318504 711590 6 vssa2
port 536 nsew ground input
rlabel metal4 s 353904 425308 354504 711590 6 vssa2
port 536 nsew ground input
rlabel metal4 s 389904 425308 390504 711590 6 vssa2
port 536 nsew ground input
rlabel metal4 s 425904 425308 426504 711590 6 vssa2
port 536 nsew ground input
rlabel metal4 s 461904 425308 462504 711590 6 vssa2
port 536 nsew ground input
rlabel metal4 s 497904 -7654 498504 711590 6 vssa2
port 536 nsew ground input
rlabel metal4 s 533904 -7654 534504 711590 6 vssa2
port 536 nsew ground input
rlabel metal4 s 569904 -7654 570504 711590 6 vssa2
port 536 nsew ground input
rlabel metal4 s 592030 -7654 592650 711590 6 vssa2
port 536 nsew ground input
rlabel metal5 s -2966 -1894 586890 -1274 8 vssd1
port 537 nsew ground input
rlabel metal5 s -2966 19876 586890 20476 6 vssd1
port 537 nsew ground input
rlabel metal5 s -2966 55876 586890 56476 6 vssd1
port 537 nsew ground input
rlabel metal5 s -2966 91876 586890 92476 6 vssd1
port 537 nsew ground input
rlabel metal5 s -2966 127876 586890 128476 6 vssd1
port 537 nsew ground input
rlabel metal5 s -2966 163876 586890 164476 6 vssd1
port 537 nsew ground input
rlabel metal5 s -2966 199876 586890 200476 6 vssd1
port 537 nsew ground input
rlabel metal5 s -2966 235876 586890 236476 6 vssd1
port 537 nsew ground input
rlabel metal5 s -2966 271876 586890 272476 6 vssd1
port 537 nsew ground input
rlabel metal5 s -2966 307876 586890 308476 6 vssd1
port 537 nsew ground input
rlabel metal5 s -2966 343876 586890 344476 6 vssd1
port 537 nsew ground input
rlabel metal5 s -2966 379876 586890 380476 6 vssd1
port 537 nsew ground input
rlabel metal5 s -2966 415876 586890 416476 6 vssd1
port 537 nsew ground input
rlabel metal5 s -2966 451876 586890 452476 6 vssd1
port 537 nsew ground input
rlabel metal5 s -2966 487876 586890 488476 6 vssd1
port 537 nsew ground input
rlabel metal5 s -2966 523876 586890 524476 6 vssd1
port 537 nsew ground input
rlabel metal5 s -2966 559876 586890 560476 6 vssd1
port 537 nsew ground input
rlabel metal5 s -2966 595876 586890 596476 6 vssd1
port 537 nsew ground input
rlabel metal5 s -2966 631876 586890 632476 6 vssd1
port 537 nsew ground input
rlabel metal5 s -2966 667876 586890 668476 6 vssd1
port 537 nsew ground input
rlabel metal5 s -2966 705210 586890 705830 6 vssd1
port 537 nsew ground input
rlabel metal4 s 54804 -1894 55404 38000 6 vssd1
port 537 nsew ground input
rlabel metal4 s 90804 -1894 91404 38000 6 vssd1
port 537 nsew ground input
rlabel metal4 s 126804 -1894 127404 38000 6 vssd1
port 537 nsew ground input
rlabel metal4 s 162804 -1894 163404 38000 6 vssd1
port 537 nsew ground input
rlabel metal4 s 198804 -1894 199404 38000 6 vssd1
port 537 nsew ground input
rlabel metal4 s 234804 -1894 235404 38000 6 vssd1
port 537 nsew ground input
rlabel metal4 s 54804 243568 55404 338000 6 vssd1
port 537 nsew ground input
rlabel metal4 s 90804 243568 91404 338000 6 vssd1
port 537 nsew ground input
rlabel metal4 s 126804 243568 127404 338000 6 vssd1
port 537 nsew ground input
rlabel metal4 s 162804 243568 163404 338000 6 vssd1
port 537 nsew ground input
rlabel metal4 s 342804 -1894 343404 338000 6 vssd1
port 537 nsew ground input
rlabel metal4 s 378804 -1894 379404 338000 6 vssd1
port 537 nsew ground input
rlabel metal4 s 414804 -1894 415404 338000 6 vssd1
port 537 nsew ground input
rlabel metal4 s 450804 -1894 451404 338000 6 vssd1
port 537 nsew ground input
rlabel metal4 s -2966 -1894 -2346 705830 4 vssd1
port 537 nsew ground input
rlabel metal4 s 18804 -1894 19404 705830 6 vssd1
port 537 nsew ground input
rlabel metal4 s 54804 425308 55404 705830 6 vssd1
port 537 nsew ground input
rlabel metal4 s 90804 425308 91404 705830 6 vssd1
port 537 nsew ground input
rlabel metal4 s 126804 425308 127404 705830 6 vssd1
port 537 nsew ground input
rlabel metal4 s 162804 425308 163404 705830 6 vssd1
port 537 nsew ground input
rlabel metal4 s 198804 243568 199404 705830 6 vssd1
port 537 nsew ground input
rlabel metal4 s 234804 243568 235404 705830 6 vssd1
port 537 nsew ground input
rlabel metal4 s 270804 -1894 271404 705830 6 vssd1
port 537 nsew ground input
rlabel metal4 s 306804 -1894 307404 705830 6 vssd1
port 537 nsew ground input
rlabel metal4 s 342804 425308 343404 705830 6 vssd1
port 537 nsew ground input
rlabel metal4 s 378804 425308 379404 705830 6 vssd1
port 537 nsew ground input
rlabel metal4 s 414804 425308 415404 705830 6 vssd1
port 537 nsew ground input
rlabel metal4 s 450804 425308 451404 705830 6 vssd1
port 537 nsew ground input
rlabel metal4 s 486804 -1894 487404 705830 6 vssd1
port 537 nsew ground input
rlabel metal4 s 522804 -1894 523404 705830 6 vssd1
port 537 nsew ground input
rlabel metal4 s 558804 -1894 559404 705830 6 vssd1
port 537 nsew ground input
rlabel metal4 s 586270 -1894 586890 705830 6 vssd1
port 537 nsew ground input
rlabel metal5 s -4886 -3814 588810 -3194 8 vssd2
port 538 nsew ground input
rlabel metal5 s -4886 23576 588810 24176 6 vssd2
port 538 nsew ground input
rlabel metal5 s -4886 59576 588810 60176 6 vssd2
port 538 nsew ground input
rlabel metal5 s -4886 95576 588810 96176 6 vssd2
port 538 nsew ground input
rlabel metal5 s -4886 131576 588810 132176 6 vssd2
port 538 nsew ground input
rlabel metal5 s -4886 167576 588810 168176 6 vssd2
port 538 nsew ground input
rlabel metal5 s -4886 203576 588810 204176 6 vssd2
port 538 nsew ground input
rlabel metal5 s -4886 239576 588810 240176 6 vssd2
port 538 nsew ground input
rlabel metal5 s -4886 275576 588810 276176 6 vssd2
port 538 nsew ground input
rlabel metal5 s -4886 311576 588810 312176 6 vssd2
port 538 nsew ground input
rlabel metal5 s -4886 347576 588810 348176 6 vssd2
port 538 nsew ground input
rlabel metal5 s -4886 383576 588810 384176 6 vssd2
port 538 nsew ground input
rlabel metal5 s -4886 419576 588810 420176 6 vssd2
port 538 nsew ground input
rlabel metal5 s -4886 455576 588810 456176 6 vssd2
port 538 nsew ground input
rlabel metal5 s -4886 491576 588810 492176 6 vssd2
port 538 nsew ground input
rlabel metal5 s -4886 527576 588810 528176 6 vssd2
port 538 nsew ground input
rlabel metal5 s -4886 563576 588810 564176 6 vssd2
port 538 nsew ground input
rlabel metal5 s -4886 599576 588810 600176 6 vssd2
port 538 nsew ground input
rlabel metal5 s -4886 635576 588810 636176 6 vssd2
port 538 nsew ground input
rlabel metal5 s -4886 671576 588810 672176 6 vssd2
port 538 nsew ground input
rlabel metal5 s -4886 707130 588810 707750 6 vssd2
port 538 nsew ground input
rlabel metal4 s 58504 -3814 59104 38000 6 vssd2
port 538 nsew ground input
rlabel metal4 s 94504 -3814 95104 38000 6 vssd2
port 538 nsew ground input
rlabel metal4 s 130504 -3814 131104 38000 6 vssd2
port 538 nsew ground input
rlabel metal4 s 166504 -3814 167104 38000 6 vssd2
port 538 nsew ground input
rlabel metal4 s 202504 -3814 203104 38000 6 vssd2
port 538 nsew ground input
rlabel metal4 s 238504 -3814 239104 38000 6 vssd2
port 538 nsew ground input
rlabel metal4 s 58504 243568 59104 338000 6 vssd2
port 538 nsew ground input
rlabel metal4 s 94504 243568 95104 338000 6 vssd2
port 538 nsew ground input
rlabel metal4 s 130504 243568 131104 338000 6 vssd2
port 538 nsew ground input
rlabel metal4 s 166504 243568 167104 338000 6 vssd2
port 538 nsew ground input
rlabel metal4 s 346504 -3814 347104 338000 6 vssd2
port 538 nsew ground input
rlabel metal4 s 382504 -3814 383104 338000 6 vssd2
port 538 nsew ground input
rlabel metal4 s 418504 -3814 419104 338000 6 vssd2
port 538 nsew ground input
rlabel metal4 s 454504 -3814 455104 338000 6 vssd2
port 538 nsew ground input
rlabel metal4 s -4886 -3814 -4266 707750 4 vssd2
port 538 nsew ground input
rlabel metal4 s 22504 -3814 23104 707750 6 vssd2
port 538 nsew ground input
rlabel metal4 s 58504 425308 59104 707750 6 vssd2
port 538 nsew ground input
rlabel metal4 s 94504 425308 95104 707750 6 vssd2
port 538 nsew ground input
rlabel metal4 s 130504 425308 131104 707750 6 vssd2
port 538 nsew ground input
rlabel metal4 s 166504 425308 167104 707750 6 vssd2
port 538 nsew ground input
rlabel metal4 s 202504 243568 203104 707750 6 vssd2
port 538 nsew ground input
rlabel metal4 s 238504 243568 239104 707750 6 vssd2
port 538 nsew ground input
rlabel metal4 s 274504 -3814 275104 707750 6 vssd2
port 538 nsew ground input
rlabel metal4 s 310504 -3814 311104 707750 6 vssd2
port 538 nsew ground input
rlabel metal4 s 346504 425308 347104 707750 6 vssd2
port 538 nsew ground input
rlabel metal4 s 382504 425308 383104 707750 6 vssd2
port 538 nsew ground input
rlabel metal4 s 418504 425308 419104 707750 6 vssd2
port 538 nsew ground input
rlabel metal4 s 454504 425308 455104 707750 6 vssd2
port 538 nsew ground input
rlabel metal4 s 490504 -3814 491104 707750 6 vssd2
port 538 nsew ground input
rlabel metal4 s 526504 -3814 527104 707750 6 vssd2
port 538 nsew ground input
rlabel metal4 s 562504 -3814 563104 707750 6 vssd2
port 538 nsew ground input
rlabel metal4 s 588190 -3814 588810 707750 6 vssd2
port 538 nsew ground input
rlabel metal2 s 542 -960 654 480 8 wb_clk_i
port 539 nsew signal input
rlabel metal2 s 1646 -960 1758 480 8 wb_rst_i
port 540 nsew signal input
rlabel metal2 s 2842 -960 2954 480 8 wbs_ack_o
port 541 nsew signal tristate
rlabel metal2 s 7626 -960 7738 480 8 wbs_adr_i[0]
port 542 nsew signal input
rlabel metal2 s 47830 -960 47942 480 8 wbs_adr_i[10]
port 543 nsew signal input
rlabel metal2 s 51326 -960 51438 480 8 wbs_adr_i[11]
port 544 nsew signal input
rlabel metal2 s 54914 -960 55026 480 8 wbs_adr_i[12]
port 545 nsew signal input
rlabel metal2 s 58410 -960 58522 480 8 wbs_adr_i[13]
port 546 nsew signal input
rlabel metal2 s 61998 -960 62110 480 8 wbs_adr_i[14]
port 547 nsew signal input
rlabel metal2 s 65494 -960 65606 480 8 wbs_adr_i[15]
port 548 nsew signal input
rlabel metal2 s 69082 -960 69194 480 8 wbs_adr_i[16]
port 549 nsew signal input
rlabel metal2 s 72578 -960 72690 480 8 wbs_adr_i[17]
port 550 nsew signal input
rlabel metal2 s 76166 -960 76278 480 8 wbs_adr_i[18]
port 551 nsew signal input
rlabel metal2 s 79662 -960 79774 480 8 wbs_adr_i[19]
port 552 nsew signal input
rlabel metal2 s 12318 -960 12430 480 8 wbs_adr_i[1]
port 553 nsew signal input
rlabel metal2 s 83250 -960 83362 480 8 wbs_adr_i[20]
port 554 nsew signal input
rlabel metal2 s 86838 -960 86950 480 8 wbs_adr_i[21]
port 555 nsew signal input
rlabel metal2 s 90334 -960 90446 480 8 wbs_adr_i[22]
port 556 nsew signal input
rlabel metal2 s 93922 -960 94034 480 8 wbs_adr_i[23]
port 557 nsew signal input
rlabel metal2 s 97418 -960 97530 480 8 wbs_adr_i[24]
port 558 nsew signal input
rlabel metal2 s 101006 -960 101118 480 8 wbs_adr_i[25]
port 559 nsew signal input
rlabel metal2 s 104502 -960 104614 480 8 wbs_adr_i[26]
port 560 nsew signal input
rlabel metal2 s 108090 -960 108202 480 8 wbs_adr_i[27]
port 561 nsew signal input
rlabel metal2 s 111586 -960 111698 480 8 wbs_adr_i[28]
port 562 nsew signal input
rlabel metal2 s 115174 -960 115286 480 8 wbs_adr_i[29]
port 563 nsew signal input
rlabel metal2 s 17010 -960 17122 480 8 wbs_adr_i[2]
port 564 nsew signal input
rlabel metal2 s 118762 -960 118874 480 8 wbs_adr_i[30]
port 565 nsew signal input
rlabel metal2 s 122258 -960 122370 480 8 wbs_adr_i[31]
port 566 nsew signal input
rlabel metal2 s 21794 -960 21906 480 8 wbs_adr_i[3]
port 567 nsew signal input
rlabel metal2 s 26486 -960 26598 480 8 wbs_adr_i[4]
port 568 nsew signal input
rlabel metal2 s 30074 -960 30186 480 8 wbs_adr_i[5]
port 569 nsew signal input
rlabel metal2 s 33570 -960 33682 480 8 wbs_adr_i[6]
port 570 nsew signal input
rlabel metal2 s 37158 -960 37270 480 8 wbs_adr_i[7]
port 571 nsew signal input
rlabel metal2 s 40654 -960 40766 480 8 wbs_adr_i[8]
port 572 nsew signal input
rlabel metal2 s 44242 -960 44354 480 8 wbs_adr_i[9]
port 573 nsew signal input
rlabel metal2 s 4038 -960 4150 480 8 wbs_cyc_i
port 574 nsew signal input
rlabel metal2 s 8730 -960 8842 480 8 wbs_dat_i[0]
port 575 nsew signal input
rlabel metal2 s 48934 -960 49046 480 8 wbs_dat_i[10]
port 576 nsew signal input
rlabel metal2 s 52522 -960 52634 480 8 wbs_dat_i[11]
port 577 nsew signal input
rlabel metal2 s 56018 -960 56130 480 8 wbs_dat_i[12]
port 578 nsew signal input
rlabel metal2 s 59606 -960 59718 480 8 wbs_dat_i[13]
port 579 nsew signal input
rlabel metal2 s 63194 -960 63306 480 8 wbs_dat_i[14]
port 580 nsew signal input
rlabel metal2 s 66690 -960 66802 480 8 wbs_dat_i[15]
port 581 nsew signal input
rlabel metal2 s 70278 -960 70390 480 8 wbs_dat_i[16]
port 582 nsew signal input
rlabel metal2 s 73774 -960 73886 480 8 wbs_dat_i[17]
port 583 nsew signal input
rlabel metal2 s 77362 -960 77474 480 8 wbs_dat_i[18]
port 584 nsew signal input
rlabel metal2 s 80858 -960 80970 480 8 wbs_dat_i[19]
port 585 nsew signal input
rlabel metal2 s 13514 -960 13626 480 8 wbs_dat_i[1]
port 586 nsew signal input
rlabel metal2 s 84446 -960 84558 480 8 wbs_dat_i[20]
port 587 nsew signal input
rlabel metal2 s 87942 -960 88054 480 8 wbs_dat_i[21]
port 588 nsew signal input
rlabel metal2 s 91530 -960 91642 480 8 wbs_dat_i[22]
port 589 nsew signal input
rlabel metal2 s 95118 -960 95230 480 8 wbs_dat_i[23]
port 590 nsew signal input
rlabel metal2 s 98614 -960 98726 480 8 wbs_dat_i[24]
port 591 nsew signal input
rlabel metal2 s 102202 -960 102314 480 8 wbs_dat_i[25]
port 592 nsew signal input
rlabel metal2 s 105698 -960 105810 480 8 wbs_dat_i[26]
port 593 nsew signal input
rlabel metal2 s 109286 -960 109398 480 8 wbs_dat_i[27]
port 594 nsew signal input
rlabel metal2 s 112782 -960 112894 480 8 wbs_dat_i[28]
port 595 nsew signal input
rlabel metal2 s 116370 -960 116482 480 8 wbs_dat_i[29]
port 596 nsew signal input
rlabel metal2 s 18206 -960 18318 480 8 wbs_dat_i[2]
port 597 nsew signal input
rlabel metal2 s 119866 -960 119978 480 8 wbs_dat_i[30]
port 598 nsew signal input
rlabel metal2 s 123454 -960 123566 480 8 wbs_dat_i[31]
port 599 nsew signal input
rlabel metal2 s 22990 -960 23102 480 8 wbs_dat_i[3]
port 600 nsew signal input
rlabel metal2 s 27682 -960 27794 480 8 wbs_dat_i[4]
port 601 nsew signal input
rlabel metal2 s 31270 -960 31382 480 8 wbs_dat_i[5]
port 602 nsew signal input
rlabel metal2 s 34766 -960 34878 480 8 wbs_dat_i[6]
port 603 nsew signal input
rlabel metal2 s 38354 -960 38466 480 8 wbs_dat_i[7]
port 604 nsew signal input
rlabel metal2 s 41850 -960 41962 480 8 wbs_dat_i[8]
port 605 nsew signal input
rlabel metal2 s 45438 -960 45550 480 8 wbs_dat_i[9]
port 606 nsew signal input
rlabel metal2 s 9926 -960 10038 480 8 wbs_dat_o[0]
port 607 nsew signal tristate
rlabel metal2 s 50130 -960 50242 480 8 wbs_dat_o[10]
port 608 nsew signal tristate
rlabel metal2 s 53718 -960 53830 480 8 wbs_dat_o[11]
port 609 nsew signal tristate
rlabel metal2 s 57214 -960 57326 480 8 wbs_dat_o[12]
port 610 nsew signal tristate
rlabel metal2 s 60802 -960 60914 480 8 wbs_dat_o[13]
port 611 nsew signal tristate
rlabel metal2 s 64298 -960 64410 480 8 wbs_dat_o[14]
port 612 nsew signal tristate
rlabel metal2 s 67886 -960 67998 480 8 wbs_dat_o[15]
port 613 nsew signal tristate
rlabel metal2 s 71474 -960 71586 480 8 wbs_dat_o[16]
port 614 nsew signal tristate
rlabel metal2 s 74970 -960 75082 480 8 wbs_dat_o[17]
port 615 nsew signal tristate
rlabel metal2 s 78558 -960 78670 480 8 wbs_dat_o[18]
port 616 nsew signal tristate
rlabel metal2 s 82054 -960 82166 480 8 wbs_dat_o[19]
port 617 nsew signal tristate
rlabel metal2 s 14710 -960 14822 480 8 wbs_dat_o[1]
port 618 nsew signal tristate
rlabel metal2 s 85642 -960 85754 480 8 wbs_dat_o[20]
port 619 nsew signal tristate
rlabel metal2 s 89138 -960 89250 480 8 wbs_dat_o[21]
port 620 nsew signal tristate
rlabel metal2 s 92726 -960 92838 480 8 wbs_dat_o[22]
port 621 nsew signal tristate
rlabel metal2 s 96222 -960 96334 480 8 wbs_dat_o[23]
port 622 nsew signal tristate
rlabel metal2 s 99810 -960 99922 480 8 wbs_dat_o[24]
port 623 nsew signal tristate
rlabel metal2 s 103306 -960 103418 480 8 wbs_dat_o[25]
port 624 nsew signal tristate
rlabel metal2 s 106894 -960 107006 480 8 wbs_dat_o[26]
port 625 nsew signal tristate
rlabel metal2 s 110482 -960 110594 480 8 wbs_dat_o[27]
port 626 nsew signal tristate
rlabel metal2 s 113978 -960 114090 480 8 wbs_dat_o[28]
port 627 nsew signal tristate
rlabel metal2 s 117566 -960 117678 480 8 wbs_dat_o[29]
port 628 nsew signal tristate
rlabel metal2 s 19402 -960 19514 480 8 wbs_dat_o[2]
port 629 nsew signal tristate
rlabel metal2 s 121062 -960 121174 480 8 wbs_dat_o[30]
port 630 nsew signal tristate
rlabel metal2 s 124650 -960 124762 480 8 wbs_dat_o[31]
port 631 nsew signal tristate
rlabel metal2 s 24186 -960 24298 480 8 wbs_dat_o[3]
port 632 nsew signal tristate
rlabel metal2 s 28878 -960 28990 480 8 wbs_dat_o[4]
port 633 nsew signal tristate
rlabel metal2 s 32374 -960 32486 480 8 wbs_dat_o[5]
port 634 nsew signal tristate
rlabel metal2 s 35962 -960 36074 480 8 wbs_dat_o[6]
port 635 nsew signal tristate
rlabel metal2 s 39550 -960 39662 480 8 wbs_dat_o[7]
port 636 nsew signal tristate
rlabel metal2 s 43046 -960 43158 480 8 wbs_dat_o[8]
port 637 nsew signal tristate
rlabel metal2 s 46634 -960 46746 480 8 wbs_dat_o[9]
port 638 nsew signal tristate
rlabel metal2 s 11122 -960 11234 480 8 wbs_sel_i[0]
port 639 nsew signal input
rlabel metal2 s 15906 -960 16018 480 8 wbs_sel_i[1]
port 640 nsew signal input
rlabel metal2 s 20598 -960 20710 480 8 wbs_sel_i[2]
port 641 nsew signal input
rlabel metal2 s 25290 -960 25402 480 8 wbs_sel_i[3]
port 642 nsew signal input
rlabel metal2 s 5234 -960 5346 480 8 wbs_stb_i
port 643 nsew signal input
rlabel metal2 s 6430 -960 6542 480 8 wbs_we_i
port 644 nsew signal input
<< properties >>
string FIXED_BBOX 0 0 584000 704000
<< end >>
