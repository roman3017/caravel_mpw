magic
tech sky130A
magscale 1 2
timestamp 1643614346
<< obsli1 >>
rect 1104 2159 197771 198033
<< obsm1 >>
rect 566 1504 197878 198280
<< metal2 >>
rect 662 199469 718 200269
rect 1950 199469 2006 200269
rect 3238 199469 3294 200269
rect 4526 199469 4582 200269
rect 5814 199469 5870 200269
rect 7102 199469 7158 200269
rect 8390 199469 8446 200269
rect 9678 199469 9734 200269
rect 10966 199469 11022 200269
rect 12254 199469 12310 200269
rect 13542 199469 13598 200269
rect 14830 199469 14886 200269
rect 16118 199469 16174 200269
rect 17498 199469 17554 200269
rect 18786 199469 18842 200269
rect 20074 199469 20130 200269
rect 21362 199469 21418 200269
rect 22650 199469 22706 200269
rect 23938 199469 23994 200269
rect 25226 199469 25282 200269
rect 26514 199469 26570 200269
rect 27802 199469 27858 200269
rect 29090 199469 29146 200269
rect 30378 199469 30434 200269
rect 31666 199469 31722 200269
rect 32954 199469 33010 200269
rect 34334 199469 34390 200269
rect 35622 199469 35678 200269
rect 36910 199469 36966 200269
rect 38198 199469 38254 200269
rect 39486 199469 39542 200269
rect 40774 199469 40830 200269
rect 42062 199469 42118 200269
rect 43350 199469 43406 200269
rect 44638 199469 44694 200269
rect 45926 199469 45982 200269
rect 47214 199469 47270 200269
rect 48502 199469 48558 200269
rect 49790 199469 49846 200269
rect 51170 199469 51226 200269
rect 52458 199469 52514 200269
rect 53746 199469 53802 200269
rect 55034 199469 55090 200269
rect 56322 199469 56378 200269
rect 57610 199469 57666 200269
rect 58898 199469 58954 200269
rect 60186 199469 60242 200269
rect 61474 199469 61530 200269
rect 62762 199469 62818 200269
rect 64050 199469 64106 200269
rect 65338 199469 65394 200269
rect 66718 199469 66774 200269
rect 68006 199469 68062 200269
rect 69294 199469 69350 200269
rect 70582 199469 70638 200269
rect 71870 199469 71926 200269
rect 73158 199469 73214 200269
rect 74446 199469 74502 200269
rect 75734 199469 75790 200269
rect 77022 199469 77078 200269
rect 78310 199469 78366 200269
rect 79598 199469 79654 200269
rect 80886 199469 80942 200269
rect 82174 199469 82230 200269
rect 83554 199469 83610 200269
rect 84842 199469 84898 200269
rect 86130 199469 86186 200269
rect 87418 199469 87474 200269
rect 88706 199469 88762 200269
rect 89994 199469 90050 200269
rect 91282 199469 91338 200269
rect 92570 199469 92626 200269
rect 93858 199469 93914 200269
rect 95146 199469 95202 200269
rect 96434 199469 96490 200269
rect 97722 199469 97778 200269
rect 99010 199469 99066 200269
rect 100390 199469 100446 200269
rect 101678 199469 101734 200269
rect 102966 199469 103022 200269
rect 104254 199469 104310 200269
rect 105542 199469 105598 200269
rect 106830 199469 106886 200269
rect 108118 199469 108174 200269
rect 109406 199469 109462 200269
rect 110694 199469 110750 200269
rect 111982 199469 112038 200269
rect 113270 199469 113326 200269
rect 114558 199469 114614 200269
rect 115846 199469 115902 200269
rect 117226 199469 117282 200269
rect 118514 199469 118570 200269
rect 119802 199469 119858 200269
rect 121090 199469 121146 200269
rect 122378 199469 122434 200269
rect 123666 199469 123722 200269
rect 124954 199469 125010 200269
rect 126242 199469 126298 200269
rect 127530 199469 127586 200269
rect 128818 199469 128874 200269
rect 130106 199469 130162 200269
rect 131394 199469 131450 200269
rect 132774 199469 132830 200269
rect 134062 199469 134118 200269
rect 135350 199469 135406 200269
rect 136638 199469 136694 200269
rect 137926 199469 137982 200269
rect 139214 199469 139270 200269
rect 140502 199469 140558 200269
rect 141790 199469 141846 200269
rect 143078 199469 143134 200269
rect 144366 199469 144422 200269
rect 145654 199469 145710 200269
rect 146942 199469 146998 200269
rect 148230 199469 148286 200269
rect 149610 199469 149666 200269
rect 150898 199469 150954 200269
rect 152186 199469 152242 200269
rect 153474 199469 153530 200269
rect 154762 199469 154818 200269
rect 156050 199469 156106 200269
rect 157338 199469 157394 200269
rect 158626 199469 158682 200269
rect 159914 199469 159970 200269
rect 161202 199469 161258 200269
rect 162490 199469 162546 200269
rect 163778 199469 163834 200269
rect 165066 199469 165122 200269
rect 166446 199469 166502 200269
rect 167734 199469 167790 200269
rect 169022 199469 169078 200269
rect 170310 199469 170366 200269
rect 171598 199469 171654 200269
rect 172886 199469 172942 200269
rect 174174 199469 174230 200269
rect 175462 199469 175518 200269
rect 176750 199469 176806 200269
rect 178038 199469 178094 200269
rect 179326 199469 179382 200269
rect 180614 199469 180670 200269
rect 181902 199469 181958 200269
rect 183282 199469 183338 200269
rect 184570 199469 184626 200269
rect 185858 199469 185914 200269
rect 187146 199469 187202 200269
rect 188434 199469 188490 200269
rect 189722 199469 189778 200269
rect 191010 199469 191066 200269
rect 192298 199469 192354 200269
rect 193586 199469 193642 200269
rect 194874 199469 194930 200269
rect 196162 199469 196218 200269
rect 197450 199469 197506 200269
rect 570 0 626 800
rect 1766 0 1822 800
rect 3054 0 3110 800
rect 4250 0 4306 800
rect 5538 0 5594 800
rect 6734 0 6790 800
rect 8022 0 8078 800
rect 9218 0 9274 800
rect 10506 0 10562 800
rect 11702 0 11758 800
rect 12990 0 13046 800
rect 14278 0 14334 800
rect 15474 0 15530 800
rect 16762 0 16818 800
rect 17958 0 18014 800
rect 19246 0 19302 800
rect 20442 0 20498 800
rect 21730 0 21786 800
rect 22926 0 22982 800
rect 24214 0 24270 800
rect 25410 0 25466 800
rect 26698 0 26754 800
rect 27986 0 28042 800
rect 29182 0 29238 800
rect 30470 0 30526 800
rect 31666 0 31722 800
rect 32954 0 33010 800
rect 34150 0 34206 800
rect 35438 0 35494 800
rect 36634 0 36690 800
rect 37922 0 37978 800
rect 39118 0 39174 800
rect 40406 0 40462 800
rect 41694 0 41750 800
rect 42890 0 42946 800
rect 44178 0 44234 800
rect 45374 0 45430 800
rect 46662 0 46718 800
rect 47858 0 47914 800
rect 49146 0 49202 800
rect 50342 0 50398 800
rect 51630 0 51686 800
rect 52826 0 52882 800
rect 54114 0 54170 800
rect 55402 0 55458 800
rect 56598 0 56654 800
rect 57886 0 57942 800
rect 59082 0 59138 800
rect 60370 0 60426 800
rect 61566 0 61622 800
rect 62854 0 62910 800
rect 64050 0 64106 800
rect 65338 0 65394 800
rect 66626 0 66682 800
rect 67822 0 67878 800
rect 69110 0 69166 800
rect 70306 0 70362 800
rect 71594 0 71650 800
rect 72790 0 72846 800
rect 74078 0 74134 800
rect 75274 0 75330 800
rect 76562 0 76618 800
rect 77758 0 77814 800
rect 79046 0 79102 800
rect 80334 0 80390 800
rect 81530 0 81586 800
rect 82818 0 82874 800
rect 84014 0 84070 800
rect 85302 0 85358 800
rect 86498 0 86554 800
rect 87786 0 87842 800
rect 88982 0 89038 800
rect 90270 0 90326 800
rect 91466 0 91522 800
rect 92754 0 92810 800
rect 94042 0 94098 800
rect 95238 0 95294 800
rect 96526 0 96582 800
rect 97722 0 97778 800
rect 99010 0 99066 800
rect 100206 0 100262 800
rect 101494 0 101550 800
rect 102690 0 102746 800
rect 103978 0 104034 800
rect 105174 0 105230 800
rect 106462 0 106518 800
rect 107750 0 107806 800
rect 108946 0 109002 800
rect 110234 0 110290 800
rect 111430 0 111486 800
rect 112718 0 112774 800
rect 113914 0 113970 800
rect 115202 0 115258 800
rect 116398 0 116454 800
rect 117686 0 117742 800
rect 118882 0 118938 800
rect 120170 0 120226 800
rect 121458 0 121514 800
rect 122654 0 122710 800
rect 123942 0 123998 800
rect 125138 0 125194 800
rect 126426 0 126482 800
rect 127622 0 127678 800
rect 128910 0 128966 800
rect 130106 0 130162 800
rect 131394 0 131450 800
rect 132682 0 132738 800
rect 133878 0 133934 800
rect 135166 0 135222 800
rect 136362 0 136418 800
rect 137650 0 137706 800
rect 138846 0 138902 800
rect 140134 0 140190 800
rect 141330 0 141386 800
rect 142618 0 142674 800
rect 143814 0 143870 800
rect 145102 0 145158 800
rect 146390 0 146446 800
rect 147586 0 147642 800
rect 148874 0 148930 800
rect 150070 0 150126 800
rect 151358 0 151414 800
rect 152554 0 152610 800
rect 153842 0 153898 800
rect 155038 0 155094 800
rect 156326 0 156382 800
rect 157522 0 157578 800
rect 158810 0 158866 800
rect 160098 0 160154 800
rect 161294 0 161350 800
rect 162582 0 162638 800
rect 163778 0 163834 800
rect 165066 0 165122 800
rect 166262 0 166318 800
rect 167550 0 167606 800
rect 168746 0 168802 800
rect 170034 0 170090 800
rect 171230 0 171286 800
rect 172518 0 172574 800
rect 173806 0 173862 800
rect 175002 0 175058 800
rect 176290 0 176346 800
rect 177486 0 177542 800
rect 178774 0 178830 800
rect 179970 0 180026 800
rect 181258 0 181314 800
rect 182454 0 182510 800
rect 183742 0 183798 800
rect 184938 0 184994 800
rect 186226 0 186282 800
rect 187514 0 187570 800
rect 188710 0 188766 800
rect 189998 0 190054 800
rect 191194 0 191250 800
rect 192482 0 192538 800
rect 193678 0 193734 800
rect 194966 0 195022 800
rect 196162 0 196218 800
rect 197450 0 197506 800
<< obsm2 >>
rect 572 199413 606 199469
rect 774 199413 1894 199469
rect 2062 199413 3182 199469
rect 3350 199413 4470 199469
rect 4638 199413 5758 199469
rect 5926 199413 7046 199469
rect 7214 199413 8334 199469
rect 8502 199413 9622 199469
rect 9790 199413 10910 199469
rect 11078 199413 12198 199469
rect 12366 199413 13486 199469
rect 13654 199413 14774 199469
rect 14942 199413 16062 199469
rect 16230 199413 17442 199469
rect 17610 199413 18730 199469
rect 18898 199413 20018 199469
rect 20186 199413 21306 199469
rect 21474 199413 22594 199469
rect 22762 199413 23882 199469
rect 24050 199413 25170 199469
rect 25338 199413 26458 199469
rect 26626 199413 27746 199469
rect 27914 199413 29034 199469
rect 29202 199413 30322 199469
rect 30490 199413 31610 199469
rect 31778 199413 32898 199469
rect 33066 199413 34278 199469
rect 34446 199413 35566 199469
rect 35734 199413 36854 199469
rect 37022 199413 38142 199469
rect 38310 199413 39430 199469
rect 39598 199413 40718 199469
rect 40886 199413 42006 199469
rect 42174 199413 43294 199469
rect 43462 199413 44582 199469
rect 44750 199413 45870 199469
rect 46038 199413 47158 199469
rect 47326 199413 48446 199469
rect 48614 199413 49734 199469
rect 49902 199413 51114 199469
rect 51282 199413 52402 199469
rect 52570 199413 53690 199469
rect 53858 199413 54978 199469
rect 55146 199413 56266 199469
rect 56434 199413 57554 199469
rect 57722 199413 58842 199469
rect 59010 199413 60130 199469
rect 60298 199413 61418 199469
rect 61586 199413 62706 199469
rect 62874 199413 63994 199469
rect 64162 199413 65282 199469
rect 65450 199413 66662 199469
rect 66830 199413 67950 199469
rect 68118 199413 69238 199469
rect 69406 199413 70526 199469
rect 70694 199413 71814 199469
rect 71982 199413 73102 199469
rect 73270 199413 74390 199469
rect 74558 199413 75678 199469
rect 75846 199413 76966 199469
rect 77134 199413 78254 199469
rect 78422 199413 79542 199469
rect 79710 199413 80830 199469
rect 80998 199413 82118 199469
rect 82286 199413 83498 199469
rect 83666 199413 84786 199469
rect 84954 199413 86074 199469
rect 86242 199413 87362 199469
rect 87530 199413 88650 199469
rect 88818 199413 89938 199469
rect 90106 199413 91226 199469
rect 91394 199413 92514 199469
rect 92682 199413 93802 199469
rect 93970 199413 95090 199469
rect 95258 199413 96378 199469
rect 96546 199413 97666 199469
rect 97834 199413 98954 199469
rect 99122 199413 100334 199469
rect 100502 199413 101622 199469
rect 101790 199413 102910 199469
rect 103078 199413 104198 199469
rect 104366 199413 105486 199469
rect 105654 199413 106774 199469
rect 106942 199413 108062 199469
rect 108230 199413 109350 199469
rect 109518 199413 110638 199469
rect 110806 199413 111926 199469
rect 112094 199413 113214 199469
rect 113382 199413 114502 199469
rect 114670 199413 115790 199469
rect 115958 199413 117170 199469
rect 117338 199413 118458 199469
rect 118626 199413 119746 199469
rect 119914 199413 121034 199469
rect 121202 199413 122322 199469
rect 122490 199413 123610 199469
rect 123778 199413 124898 199469
rect 125066 199413 126186 199469
rect 126354 199413 127474 199469
rect 127642 199413 128762 199469
rect 128930 199413 130050 199469
rect 130218 199413 131338 199469
rect 131506 199413 132718 199469
rect 132886 199413 134006 199469
rect 134174 199413 135294 199469
rect 135462 199413 136582 199469
rect 136750 199413 137870 199469
rect 138038 199413 139158 199469
rect 139326 199413 140446 199469
rect 140614 199413 141734 199469
rect 141902 199413 143022 199469
rect 143190 199413 144310 199469
rect 144478 199413 145598 199469
rect 145766 199413 146886 199469
rect 147054 199413 148174 199469
rect 148342 199413 149554 199469
rect 149722 199413 150842 199469
rect 151010 199413 152130 199469
rect 152298 199413 153418 199469
rect 153586 199413 154706 199469
rect 154874 199413 155994 199469
rect 156162 199413 157282 199469
rect 157450 199413 158570 199469
rect 158738 199413 159858 199469
rect 160026 199413 161146 199469
rect 161314 199413 162434 199469
rect 162602 199413 163722 199469
rect 163890 199413 165010 199469
rect 165178 199413 166390 199469
rect 166558 199413 167678 199469
rect 167846 199413 168966 199469
rect 169134 199413 170254 199469
rect 170422 199413 171542 199469
rect 171710 199413 172830 199469
rect 172998 199413 174118 199469
rect 174286 199413 175406 199469
rect 175574 199413 176694 199469
rect 176862 199413 177982 199469
rect 178150 199413 179270 199469
rect 179438 199413 180558 199469
rect 180726 199413 181846 199469
rect 182014 199413 183226 199469
rect 183394 199413 184514 199469
rect 184682 199413 185802 199469
rect 185970 199413 187090 199469
rect 187258 199413 188378 199469
rect 188546 199413 189666 199469
rect 189834 199413 190954 199469
rect 191122 199413 192242 199469
rect 192410 199413 193530 199469
rect 193698 199413 194818 199469
rect 194986 199413 196106 199469
rect 196274 199413 197394 199469
rect 197562 199413 197872 199469
rect 572 856 197872 199413
rect 682 734 1710 856
rect 1878 734 2998 856
rect 3166 734 4194 856
rect 4362 734 5482 856
rect 5650 734 6678 856
rect 6846 734 7966 856
rect 8134 734 9162 856
rect 9330 734 10450 856
rect 10618 734 11646 856
rect 11814 734 12934 856
rect 13102 734 14222 856
rect 14390 734 15418 856
rect 15586 734 16706 856
rect 16874 734 17902 856
rect 18070 734 19190 856
rect 19358 734 20386 856
rect 20554 734 21674 856
rect 21842 734 22870 856
rect 23038 734 24158 856
rect 24326 734 25354 856
rect 25522 734 26642 856
rect 26810 734 27930 856
rect 28098 734 29126 856
rect 29294 734 30414 856
rect 30582 734 31610 856
rect 31778 734 32898 856
rect 33066 734 34094 856
rect 34262 734 35382 856
rect 35550 734 36578 856
rect 36746 734 37866 856
rect 38034 734 39062 856
rect 39230 734 40350 856
rect 40518 734 41638 856
rect 41806 734 42834 856
rect 43002 734 44122 856
rect 44290 734 45318 856
rect 45486 734 46606 856
rect 46774 734 47802 856
rect 47970 734 49090 856
rect 49258 734 50286 856
rect 50454 734 51574 856
rect 51742 734 52770 856
rect 52938 734 54058 856
rect 54226 734 55346 856
rect 55514 734 56542 856
rect 56710 734 57830 856
rect 57998 734 59026 856
rect 59194 734 60314 856
rect 60482 734 61510 856
rect 61678 734 62798 856
rect 62966 734 63994 856
rect 64162 734 65282 856
rect 65450 734 66570 856
rect 66738 734 67766 856
rect 67934 734 69054 856
rect 69222 734 70250 856
rect 70418 734 71538 856
rect 71706 734 72734 856
rect 72902 734 74022 856
rect 74190 734 75218 856
rect 75386 734 76506 856
rect 76674 734 77702 856
rect 77870 734 78990 856
rect 79158 734 80278 856
rect 80446 734 81474 856
rect 81642 734 82762 856
rect 82930 734 83958 856
rect 84126 734 85246 856
rect 85414 734 86442 856
rect 86610 734 87730 856
rect 87898 734 88926 856
rect 89094 734 90214 856
rect 90382 734 91410 856
rect 91578 734 92698 856
rect 92866 734 93986 856
rect 94154 734 95182 856
rect 95350 734 96470 856
rect 96638 734 97666 856
rect 97834 734 98954 856
rect 99122 734 100150 856
rect 100318 734 101438 856
rect 101606 734 102634 856
rect 102802 734 103922 856
rect 104090 734 105118 856
rect 105286 734 106406 856
rect 106574 734 107694 856
rect 107862 734 108890 856
rect 109058 734 110178 856
rect 110346 734 111374 856
rect 111542 734 112662 856
rect 112830 734 113858 856
rect 114026 734 115146 856
rect 115314 734 116342 856
rect 116510 734 117630 856
rect 117798 734 118826 856
rect 118994 734 120114 856
rect 120282 734 121402 856
rect 121570 734 122598 856
rect 122766 734 123886 856
rect 124054 734 125082 856
rect 125250 734 126370 856
rect 126538 734 127566 856
rect 127734 734 128854 856
rect 129022 734 130050 856
rect 130218 734 131338 856
rect 131506 734 132626 856
rect 132794 734 133822 856
rect 133990 734 135110 856
rect 135278 734 136306 856
rect 136474 734 137594 856
rect 137762 734 138790 856
rect 138958 734 140078 856
rect 140246 734 141274 856
rect 141442 734 142562 856
rect 142730 734 143758 856
rect 143926 734 145046 856
rect 145214 734 146334 856
rect 146502 734 147530 856
rect 147698 734 148818 856
rect 148986 734 150014 856
rect 150182 734 151302 856
rect 151470 734 152498 856
rect 152666 734 153786 856
rect 153954 734 154982 856
rect 155150 734 156270 856
rect 156438 734 157466 856
rect 157634 734 158754 856
rect 158922 734 160042 856
rect 160210 734 161238 856
rect 161406 734 162526 856
rect 162694 734 163722 856
rect 163890 734 165010 856
rect 165178 734 166206 856
rect 166374 734 167494 856
rect 167662 734 168690 856
rect 168858 734 169978 856
rect 170146 734 171174 856
rect 171342 734 172462 856
rect 172630 734 173750 856
rect 173918 734 174946 856
rect 175114 734 176234 856
rect 176402 734 177430 856
rect 177598 734 178718 856
rect 178886 734 179914 856
rect 180082 734 181202 856
rect 181370 734 182398 856
rect 182566 734 183686 856
rect 183854 734 184882 856
rect 185050 734 186170 856
rect 186338 734 187458 856
rect 187626 734 188654 856
rect 188822 734 189942 856
rect 190110 734 191138 856
rect 191306 734 192426 856
rect 192594 734 193622 856
rect 193790 734 194910 856
rect 195078 734 196106 856
rect 196274 734 197394 856
rect 197562 734 197872 856
<< metal3 >>
rect 0 197480 800 197600
rect 197325 197208 198125 197328
rect 0 192040 800 192160
rect 197325 191360 198125 191480
rect 0 186600 800 186720
rect 197325 185512 198125 185632
rect 0 181160 800 181280
rect 197325 179528 198125 179648
rect 0 175720 800 175840
rect 197325 173680 198125 173800
rect 0 170416 800 170536
rect 197325 167832 198125 167952
rect 0 164976 800 165096
rect 197325 161848 198125 161968
rect 0 159536 800 159656
rect 197325 156000 198125 156120
rect 0 154096 800 154216
rect 197325 150152 198125 150272
rect 0 148656 800 148776
rect 197325 144168 198125 144288
rect 0 143352 800 143472
rect 197325 138320 198125 138440
rect 0 137912 800 138032
rect 0 132472 800 132592
rect 197325 132472 198125 132592
rect 0 127032 800 127152
rect 197325 126488 198125 126608
rect 0 121592 800 121712
rect 197325 120640 198125 120760
rect 0 116288 800 116408
rect 197325 114792 198125 114912
rect 0 110848 800 110968
rect 197325 108808 198125 108928
rect 0 105408 800 105528
rect 197325 102960 198125 103080
rect 0 99968 800 100088
rect 197325 97112 198125 97232
rect 0 94528 800 94648
rect 197325 91128 198125 91248
rect 0 89088 800 89208
rect 197325 85280 198125 85400
rect 0 83784 800 83904
rect 197325 79432 198125 79552
rect 0 78344 800 78464
rect 197325 73448 198125 73568
rect 0 72904 800 73024
rect 0 67464 800 67584
rect 197325 67600 198125 67720
rect 0 62024 800 62144
rect 197325 61752 198125 61872
rect 0 56720 800 56840
rect 197325 55768 198125 55888
rect 0 51280 800 51400
rect 197325 49920 198125 50040
rect 0 45840 800 45960
rect 197325 44072 198125 44192
rect 0 40400 800 40520
rect 197325 38088 198125 38208
rect 0 34960 800 35080
rect 197325 32240 198125 32360
rect 0 29656 800 29776
rect 197325 26392 198125 26512
rect 0 24216 800 24336
rect 197325 20408 198125 20528
rect 0 18776 800 18896
rect 197325 14560 198125 14680
rect 0 13336 800 13456
rect 197325 8712 198125 8832
rect 0 7896 800 8016
rect 197325 2864 198125 2984
rect 0 2592 800 2712
<< obsm3 >>
rect 800 197680 197787 198253
rect 880 197408 197787 197680
rect 880 197400 197245 197408
rect 800 197128 197245 197400
rect 800 192240 197787 197128
rect 880 191960 197787 192240
rect 800 191560 197787 191960
rect 800 191280 197245 191560
rect 800 186800 197787 191280
rect 880 186520 197787 186800
rect 800 185712 197787 186520
rect 800 185432 197245 185712
rect 800 181360 197787 185432
rect 880 181080 197787 181360
rect 800 179728 197787 181080
rect 800 179448 197245 179728
rect 800 175920 197787 179448
rect 880 175640 197787 175920
rect 800 173880 197787 175640
rect 800 173600 197245 173880
rect 800 170616 197787 173600
rect 880 170336 197787 170616
rect 800 168032 197787 170336
rect 800 167752 197245 168032
rect 800 165176 197787 167752
rect 880 164896 197787 165176
rect 800 162048 197787 164896
rect 800 161768 197245 162048
rect 800 159736 197787 161768
rect 880 159456 197787 159736
rect 800 156200 197787 159456
rect 800 155920 197245 156200
rect 800 154296 197787 155920
rect 880 154016 197787 154296
rect 800 150352 197787 154016
rect 800 150072 197245 150352
rect 800 148856 197787 150072
rect 880 148576 197787 148856
rect 800 144368 197787 148576
rect 800 144088 197245 144368
rect 800 143552 197787 144088
rect 880 143272 197787 143552
rect 800 138520 197787 143272
rect 800 138240 197245 138520
rect 800 138112 197787 138240
rect 880 137832 197787 138112
rect 800 132672 197787 137832
rect 880 132392 197245 132672
rect 800 127232 197787 132392
rect 880 126952 197787 127232
rect 800 126688 197787 126952
rect 800 126408 197245 126688
rect 800 121792 197787 126408
rect 880 121512 197787 121792
rect 800 120840 197787 121512
rect 800 120560 197245 120840
rect 800 116488 197787 120560
rect 880 116208 197787 116488
rect 800 114992 197787 116208
rect 800 114712 197245 114992
rect 800 111048 197787 114712
rect 880 110768 197787 111048
rect 800 109008 197787 110768
rect 800 108728 197245 109008
rect 800 105608 197787 108728
rect 880 105328 197787 105608
rect 800 103160 197787 105328
rect 800 102880 197245 103160
rect 800 100168 197787 102880
rect 880 99888 197787 100168
rect 800 97312 197787 99888
rect 800 97032 197245 97312
rect 800 94728 197787 97032
rect 880 94448 197787 94728
rect 800 91328 197787 94448
rect 800 91048 197245 91328
rect 800 89288 197787 91048
rect 880 89008 197787 89288
rect 800 85480 197787 89008
rect 800 85200 197245 85480
rect 800 83984 197787 85200
rect 880 83704 197787 83984
rect 800 79632 197787 83704
rect 800 79352 197245 79632
rect 800 78544 197787 79352
rect 880 78264 197787 78544
rect 800 73648 197787 78264
rect 800 73368 197245 73648
rect 800 73104 197787 73368
rect 880 72824 197787 73104
rect 800 67800 197787 72824
rect 800 67664 197245 67800
rect 880 67520 197245 67664
rect 880 67384 197787 67520
rect 800 62224 197787 67384
rect 880 61952 197787 62224
rect 880 61944 197245 61952
rect 800 61672 197245 61944
rect 800 56920 197787 61672
rect 880 56640 197787 56920
rect 800 55968 197787 56640
rect 800 55688 197245 55968
rect 800 51480 197787 55688
rect 880 51200 197787 51480
rect 800 50120 197787 51200
rect 800 49840 197245 50120
rect 800 46040 197787 49840
rect 880 45760 197787 46040
rect 800 44272 197787 45760
rect 800 43992 197245 44272
rect 800 40600 197787 43992
rect 880 40320 197787 40600
rect 800 38288 197787 40320
rect 800 38008 197245 38288
rect 800 35160 197787 38008
rect 880 34880 197787 35160
rect 800 32440 197787 34880
rect 800 32160 197245 32440
rect 800 29856 197787 32160
rect 880 29576 197787 29856
rect 800 26592 197787 29576
rect 800 26312 197245 26592
rect 800 24416 197787 26312
rect 880 24136 197787 24416
rect 800 20608 197787 24136
rect 800 20328 197245 20608
rect 800 18976 197787 20328
rect 880 18696 197787 18976
rect 800 14760 197787 18696
rect 800 14480 197245 14760
rect 800 13536 197787 14480
rect 880 13256 197787 13536
rect 800 8912 197787 13256
rect 800 8632 197245 8912
rect 800 8096 197787 8632
rect 880 7816 197787 8096
rect 800 3064 197787 7816
rect 800 2792 197245 3064
rect 880 2784 197245 2792
rect 880 2512 197787 2784
rect 800 2143 197787 2512
<< metal4 >>
rect 4208 2128 4528 198064
rect 19568 2128 19888 198064
rect 34928 2128 35248 198064
rect 50288 2128 50608 198064
rect 65648 2128 65968 198064
rect 81008 2128 81328 198064
rect 96368 2128 96688 198064
rect 111728 2128 112048 198064
rect 127088 2128 127408 198064
rect 142448 2128 142768 198064
rect 157808 2128 158128 198064
rect 173168 2128 173488 198064
rect 188528 2128 188848 198064
<< obsm4 >>
rect 21035 198144 191853 198253
rect 21035 3163 34848 198144
rect 35328 3163 50208 198144
rect 50688 3163 65568 198144
rect 66048 3163 80928 198144
rect 81408 3163 96288 198144
rect 96768 3163 111648 198144
rect 112128 3163 127008 198144
rect 127488 3163 142368 198144
rect 142848 3163 157728 198144
rect 158208 3163 173088 198144
rect 173568 3163 188448 198144
rect 188928 3163 191853 198144
<< labels >>
rlabel metal2 s 148230 199469 148286 200269 6 clk_i
port 1 nsew signal input
rlabel metal3 s 197325 2864 198125 2984 6 i_dout0[0]
port 2 nsew signal input
rlabel metal2 s 174174 199469 174230 200269 6 i_dout0[10]
port 3 nsew signal input
rlabel metal3 s 197325 91128 198125 91248 6 i_dout0[11]
port 4 nsew signal input
rlabel metal2 s 175462 199469 175518 200269 6 i_dout0[12]
port 5 nsew signal input
rlabel metal2 s 167550 0 167606 800 6 i_dout0[13]
port 6 nsew signal input
rlabel metal3 s 0 121592 800 121712 6 i_dout0[14]
port 7 nsew signal input
rlabel metal2 s 171230 0 171286 800 6 i_dout0[15]
port 8 nsew signal input
rlabel metal2 s 179326 199469 179382 200269 6 i_dout0[16]
port 9 nsew signal input
rlabel metal3 s 197325 108808 198125 108928 6 i_dout0[17]
port 10 nsew signal input
rlabel metal3 s 197325 126488 198125 126608 6 i_dout0[18]
port 11 nsew signal input
rlabel metal2 s 176290 0 176346 800 6 i_dout0[19]
port 12 nsew signal input
rlabel metal2 s 153474 199469 153530 200269 6 i_dout0[1]
port 13 nsew signal input
rlabel metal2 s 178774 0 178830 800 6 i_dout0[20]
port 14 nsew signal input
rlabel metal3 s 0 148656 800 148776 6 i_dout0[21]
port 15 nsew signal input
rlabel metal3 s 0 154096 800 154216 6 i_dout0[22]
port 16 nsew signal input
rlabel metal3 s 197325 161848 198125 161968 6 i_dout0[23]
port 17 nsew signal input
rlabel metal3 s 0 164976 800 165096 6 i_dout0[24]
port 18 nsew signal input
rlabel metal3 s 0 170416 800 170536 6 i_dout0[25]
port 19 nsew signal input
rlabel metal3 s 0 175720 800 175840 6 i_dout0[26]
port 20 nsew signal input
rlabel metal3 s 0 181160 800 181280 6 i_dout0[27]
port 21 nsew signal input
rlabel metal2 s 192482 0 192538 800 6 i_dout0[28]
port 22 nsew signal input
rlabel metal2 s 196162 199469 196218 200269 6 i_dout0[29]
port 23 nsew signal input
rlabel metal2 s 143814 0 143870 800 6 i_dout0[2]
port 24 nsew signal input
rlabel metal2 s 196162 0 196218 800 6 i_dout0[30]
port 25 nsew signal input
rlabel metal3 s 197325 191360 198125 191480 6 i_dout0[31]
port 26 nsew signal input
rlabel metal3 s 197325 38088 198125 38208 6 i_dout0[3]
port 27 nsew signal input
rlabel metal3 s 197325 49920 198125 50040 6 i_dout0[4]
port 28 nsew signal input
rlabel metal2 s 150070 0 150126 800 6 i_dout0[5]
port 29 nsew signal input
rlabel metal3 s 0 67464 800 67584 6 i_dout0[6]
port 30 nsew signal input
rlabel metal2 s 157522 0 157578 800 6 i_dout0[7]
port 31 nsew signal input
rlabel metal2 s 158810 0 158866 800 6 i_dout0[8]
port 32 nsew signal input
rlabel metal3 s 197325 73448 198125 73568 6 i_dout0[9]
port 33 nsew signal input
rlabel metal2 s 136362 0 136418 800 6 i_dout0_1[0]
port 34 nsew signal input
rlabel metal2 s 172886 199469 172942 200269 6 i_dout0_1[10]
port 35 nsew signal input
rlabel metal3 s 197325 85280 198125 85400 6 i_dout0_1[11]
port 36 nsew signal input
rlabel metal2 s 163778 0 163834 800 6 i_dout0_1[12]
port 37 nsew signal input
rlabel metal3 s 0 116288 800 116408 6 i_dout0_1[13]
port 38 nsew signal input
rlabel metal2 s 176750 199469 176806 200269 6 i_dout0_1[14]
port 39 nsew signal input
rlabel metal2 s 178038 199469 178094 200269 6 i_dout0_1[15]
port 40 nsew signal input
rlabel metal3 s 197325 102960 198125 103080 6 i_dout0_1[16]
port 41 nsew signal input
rlabel metal2 s 183282 199469 183338 200269 6 i_dout0_1[17]
port 42 nsew signal input
rlabel metal3 s 197325 120640 198125 120760 6 i_dout0_1[18]
port 43 nsew signal input
rlabel metal3 s 197325 132472 198125 132592 6 i_dout0_1[19]
port 44 nsew signal input
rlabel metal3 s 197325 20408 198125 20528 6 i_dout0_1[1]
port 45 nsew signal input
rlabel metal2 s 177486 0 177542 800 6 i_dout0_1[20]
port 46 nsew signal input
rlabel metal3 s 197325 144168 198125 144288 6 i_dout0_1[21]
port 47 nsew signal input
rlabel metal2 s 182454 0 182510 800 6 i_dout0_1[22]
port 48 nsew signal input
rlabel metal2 s 187146 199469 187202 200269 6 i_dout0_1[23]
port 49 nsew signal input
rlabel metal3 s 0 159536 800 159656 6 i_dout0_1[24]
port 50 nsew signal input
rlabel metal2 s 191010 199469 191066 200269 6 i_dout0_1[25]
port 51 nsew signal input
rlabel metal2 s 192298 199469 192354 200269 6 i_dout0_1[26]
port 52 nsew signal input
rlabel metal2 s 189998 0 190054 800 6 i_dout0_1[27]
port 53 nsew signal input
rlabel metal2 s 191194 0 191250 800 6 i_dout0_1[28]
port 54 nsew signal input
rlabel metal2 s 194874 199469 194930 200269 6 i_dout0_1[29]
port 55 nsew signal input
rlabel metal2 s 142618 0 142674 800 6 i_dout0_1[2]
port 56 nsew signal input
rlabel metal3 s 197325 185512 198125 185632 6 i_dout0_1[30]
port 57 nsew signal input
rlabel metal3 s 0 197480 800 197600 6 i_dout0_1[31]
port 58 nsew signal input
rlabel metal2 s 158626 199469 158682 200269 6 i_dout0_1[3]
port 59 nsew signal input
rlabel metal3 s 0 51280 800 51400 6 i_dout0_1[4]
port 60 nsew signal input
rlabel metal2 s 148874 0 148930 800 6 i_dout0_1[5]
port 61 nsew signal input
rlabel metal2 s 152554 0 152610 800 6 i_dout0_1[6]
port 62 nsew signal input
rlabel metal3 s 0 72904 800 73024 6 i_dout0_1[7]
port 63 nsew signal input
rlabel metal2 s 170310 199469 170366 200269 6 i_dout0_1[8]
port 64 nsew signal input
rlabel metal2 s 171598 199469 171654 200269 6 i_dout0_1[9]
port 65 nsew signal input
rlabel metal2 s 662 199469 718 200269 6 io_in[0]
port 66 nsew signal input
rlabel metal2 s 39486 199469 39542 200269 6 io_in[10]
port 67 nsew signal input
rlabel metal2 s 43350 199469 43406 200269 6 io_in[11]
port 68 nsew signal input
rlabel metal2 s 47214 199469 47270 200269 6 io_in[12]
port 69 nsew signal input
rlabel metal2 s 51170 199469 51226 200269 6 io_in[13]
port 70 nsew signal input
rlabel metal2 s 55034 199469 55090 200269 6 io_in[14]
port 71 nsew signal input
rlabel metal2 s 58898 199469 58954 200269 6 io_in[15]
port 72 nsew signal input
rlabel metal2 s 62762 199469 62818 200269 6 io_in[16]
port 73 nsew signal input
rlabel metal2 s 66718 199469 66774 200269 6 io_in[17]
port 74 nsew signal input
rlabel metal2 s 70582 199469 70638 200269 6 io_in[18]
port 75 nsew signal input
rlabel metal2 s 74446 199469 74502 200269 6 io_in[19]
port 76 nsew signal input
rlabel metal2 s 4526 199469 4582 200269 6 io_in[1]
port 77 nsew signal input
rlabel metal2 s 78310 199469 78366 200269 6 io_in[20]
port 78 nsew signal input
rlabel metal2 s 82174 199469 82230 200269 6 io_in[21]
port 79 nsew signal input
rlabel metal2 s 86130 199469 86186 200269 6 io_in[22]
port 80 nsew signal input
rlabel metal2 s 89994 199469 90050 200269 6 io_in[23]
port 81 nsew signal input
rlabel metal2 s 93858 199469 93914 200269 6 io_in[24]
port 82 nsew signal input
rlabel metal2 s 97722 199469 97778 200269 6 io_in[25]
port 83 nsew signal input
rlabel metal2 s 101678 199469 101734 200269 6 io_in[26]
port 84 nsew signal input
rlabel metal2 s 105542 199469 105598 200269 6 io_in[27]
port 85 nsew signal input
rlabel metal2 s 109406 199469 109462 200269 6 io_in[28]
port 86 nsew signal input
rlabel metal2 s 113270 199469 113326 200269 6 io_in[29]
port 87 nsew signal input
rlabel metal2 s 8390 199469 8446 200269 6 io_in[2]
port 88 nsew signal input
rlabel metal2 s 117226 199469 117282 200269 6 io_in[30]
port 89 nsew signal input
rlabel metal2 s 121090 199469 121146 200269 6 io_in[31]
port 90 nsew signal input
rlabel metal2 s 124954 199469 125010 200269 6 io_in[32]
port 91 nsew signal input
rlabel metal2 s 128818 199469 128874 200269 6 io_in[33]
port 92 nsew signal input
rlabel metal2 s 132774 199469 132830 200269 6 io_in[34]
port 93 nsew signal input
rlabel metal2 s 136638 199469 136694 200269 6 io_in[35]
port 94 nsew signal input
rlabel metal2 s 140502 199469 140558 200269 6 io_in[36]
port 95 nsew signal input
rlabel metal2 s 144366 199469 144422 200269 6 io_in[37]
port 96 nsew signal input
rlabel metal2 s 12254 199469 12310 200269 6 io_in[3]
port 97 nsew signal input
rlabel metal2 s 16118 199469 16174 200269 6 io_in[4]
port 98 nsew signal input
rlabel metal2 s 20074 199469 20130 200269 6 io_in[5]
port 99 nsew signal input
rlabel metal2 s 23938 199469 23994 200269 6 io_in[6]
port 100 nsew signal input
rlabel metal2 s 27802 199469 27858 200269 6 io_in[7]
port 101 nsew signal input
rlabel metal2 s 31666 199469 31722 200269 6 io_in[8]
port 102 nsew signal input
rlabel metal2 s 35622 199469 35678 200269 6 io_in[9]
port 103 nsew signal input
rlabel metal2 s 1950 199469 2006 200269 6 io_oeb[0]
port 104 nsew signal output
rlabel metal2 s 40774 199469 40830 200269 6 io_oeb[10]
port 105 nsew signal output
rlabel metal2 s 44638 199469 44694 200269 6 io_oeb[11]
port 106 nsew signal output
rlabel metal2 s 48502 199469 48558 200269 6 io_oeb[12]
port 107 nsew signal output
rlabel metal2 s 52458 199469 52514 200269 6 io_oeb[13]
port 108 nsew signal output
rlabel metal2 s 56322 199469 56378 200269 6 io_oeb[14]
port 109 nsew signal output
rlabel metal2 s 60186 199469 60242 200269 6 io_oeb[15]
port 110 nsew signal output
rlabel metal2 s 64050 199469 64106 200269 6 io_oeb[16]
port 111 nsew signal output
rlabel metal2 s 68006 199469 68062 200269 6 io_oeb[17]
port 112 nsew signal output
rlabel metal2 s 71870 199469 71926 200269 6 io_oeb[18]
port 113 nsew signal output
rlabel metal2 s 75734 199469 75790 200269 6 io_oeb[19]
port 114 nsew signal output
rlabel metal2 s 5814 199469 5870 200269 6 io_oeb[1]
port 115 nsew signal output
rlabel metal2 s 79598 199469 79654 200269 6 io_oeb[20]
port 116 nsew signal output
rlabel metal2 s 83554 199469 83610 200269 6 io_oeb[21]
port 117 nsew signal output
rlabel metal2 s 87418 199469 87474 200269 6 io_oeb[22]
port 118 nsew signal output
rlabel metal2 s 91282 199469 91338 200269 6 io_oeb[23]
port 119 nsew signal output
rlabel metal2 s 95146 199469 95202 200269 6 io_oeb[24]
port 120 nsew signal output
rlabel metal2 s 99010 199469 99066 200269 6 io_oeb[25]
port 121 nsew signal output
rlabel metal2 s 102966 199469 103022 200269 6 io_oeb[26]
port 122 nsew signal output
rlabel metal2 s 106830 199469 106886 200269 6 io_oeb[27]
port 123 nsew signal output
rlabel metal2 s 110694 199469 110750 200269 6 io_oeb[28]
port 124 nsew signal output
rlabel metal2 s 114558 199469 114614 200269 6 io_oeb[29]
port 125 nsew signal output
rlabel metal2 s 9678 199469 9734 200269 6 io_oeb[2]
port 126 nsew signal output
rlabel metal2 s 118514 199469 118570 200269 6 io_oeb[30]
port 127 nsew signal output
rlabel metal2 s 122378 199469 122434 200269 6 io_oeb[31]
port 128 nsew signal output
rlabel metal2 s 126242 199469 126298 200269 6 io_oeb[32]
port 129 nsew signal output
rlabel metal2 s 130106 199469 130162 200269 6 io_oeb[33]
port 130 nsew signal output
rlabel metal2 s 134062 199469 134118 200269 6 io_oeb[34]
port 131 nsew signal output
rlabel metal2 s 137926 199469 137982 200269 6 io_oeb[35]
port 132 nsew signal output
rlabel metal2 s 141790 199469 141846 200269 6 io_oeb[36]
port 133 nsew signal output
rlabel metal2 s 145654 199469 145710 200269 6 io_oeb[37]
port 134 nsew signal output
rlabel metal2 s 13542 199469 13598 200269 6 io_oeb[3]
port 135 nsew signal output
rlabel metal2 s 17498 199469 17554 200269 6 io_oeb[4]
port 136 nsew signal output
rlabel metal2 s 21362 199469 21418 200269 6 io_oeb[5]
port 137 nsew signal output
rlabel metal2 s 25226 199469 25282 200269 6 io_oeb[6]
port 138 nsew signal output
rlabel metal2 s 29090 199469 29146 200269 6 io_oeb[7]
port 139 nsew signal output
rlabel metal2 s 32954 199469 33010 200269 6 io_oeb[8]
port 140 nsew signal output
rlabel metal2 s 36910 199469 36966 200269 6 io_oeb[9]
port 141 nsew signal output
rlabel metal2 s 3238 199469 3294 200269 6 io_out[0]
port 142 nsew signal output
rlabel metal2 s 42062 199469 42118 200269 6 io_out[10]
port 143 nsew signal output
rlabel metal2 s 45926 199469 45982 200269 6 io_out[11]
port 144 nsew signal output
rlabel metal2 s 49790 199469 49846 200269 6 io_out[12]
port 145 nsew signal output
rlabel metal2 s 53746 199469 53802 200269 6 io_out[13]
port 146 nsew signal output
rlabel metal2 s 57610 199469 57666 200269 6 io_out[14]
port 147 nsew signal output
rlabel metal2 s 61474 199469 61530 200269 6 io_out[15]
port 148 nsew signal output
rlabel metal2 s 65338 199469 65394 200269 6 io_out[16]
port 149 nsew signal output
rlabel metal2 s 69294 199469 69350 200269 6 io_out[17]
port 150 nsew signal output
rlabel metal2 s 73158 199469 73214 200269 6 io_out[18]
port 151 nsew signal output
rlabel metal2 s 77022 199469 77078 200269 6 io_out[19]
port 152 nsew signal output
rlabel metal2 s 7102 199469 7158 200269 6 io_out[1]
port 153 nsew signal output
rlabel metal2 s 80886 199469 80942 200269 6 io_out[20]
port 154 nsew signal output
rlabel metal2 s 84842 199469 84898 200269 6 io_out[21]
port 155 nsew signal output
rlabel metal2 s 88706 199469 88762 200269 6 io_out[22]
port 156 nsew signal output
rlabel metal2 s 92570 199469 92626 200269 6 io_out[23]
port 157 nsew signal output
rlabel metal2 s 96434 199469 96490 200269 6 io_out[24]
port 158 nsew signal output
rlabel metal2 s 100390 199469 100446 200269 6 io_out[25]
port 159 nsew signal output
rlabel metal2 s 104254 199469 104310 200269 6 io_out[26]
port 160 nsew signal output
rlabel metal2 s 108118 199469 108174 200269 6 io_out[27]
port 161 nsew signal output
rlabel metal2 s 111982 199469 112038 200269 6 io_out[28]
port 162 nsew signal output
rlabel metal2 s 115846 199469 115902 200269 6 io_out[29]
port 163 nsew signal output
rlabel metal2 s 10966 199469 11022 200269 6 io_out[2]
port 164 nsew signal output
rlabel metal2 s 119802 199469 119858 200269 6 io_out[30]
port 165 nsew signal output
rlabel metal2 s 123666 199469 123722 200269 6 io_out[31]
port 166 nsew signal output
rlabel metal2 s 127530 199469 127586 200269 6 io_out[32]
port 167 nsew signal output
rlabel metal2 s 131394 199469 131450 200269 6 io_out[33]
port 168 nsew signal output
rlabel metal2 s 135350 199469 135406 200269 6 io_out[34]
port 169 nsew signal output
rlabel metal2 s 139214 199469 139270 200269 6 io_out[35]
port 170 nsew signal output
rlabel metal2 s 143078 199469 143134 200269 6 io_out[36]
port 171 nsew signal output
rlabel metal2 s 146942 199469 146998 200269 6 io_out[37]
port 172 nsew signal output
rlabel metal2 s 14830 199469 14886 200269 6 io_out[3]
port 173 nsew signal output
rlabel metal2 s 18786 199469 18842 200269 6 io_out[4]
port 174 nsew signal output
rlabel metal2 s 22650 199469 22706 200269 6 io_out[5]
port 175 nsew signal output
rlabel metal2 s 26514 199469 26570 200269 6 io_out[6]
port 176 nsew signal output
rlabel metal2 s 30378 199469 30434 200269 6 io_out[7]
port 177 nsew signal output
rlabel metal2 s 34334 199469 34390 200269 6 io_out[8]
port 178 nsew signal output
rlabel metal2 s 38198 199469 38254 200269 6 io_out[9]
port 179 nsew signal output
rlabel metal2 s 132682 0 132738 800 6 irq[0]
port 180 nsew signal output
rlabel metal2 s 133878 0 133934 800 6 irq[1]
port 181 nsew signal output
rlabel metal2 s 135166 0 135222 800 6 irq[2]
port 182 nsew signal output
rlabel metal3 s 0 2592 800 2712 6 o_csb0
port 183 nsew signal output
rlabel metal3 s 0 7896 800 8016 6 o_csb0_1
port 184 nsew signal output
rlabel metal2 s 137650 0 137706 800 6 o_din0[0]
port 185 nsew signal output
rlabel metal3 s 0 105408 800 105528 6 o_din0[10]
port 186 nsew signal output
rlabel metal2 s 162582 0 162638 800 6 o_din0[11]
port 187 nsew signal output
rlabel metal2 s 166262 0 166318 800 6 o_din0[12]
port 188 nsew signal output
rlabel metal2 s 170034 0 170090 800 6 o_din0[13]
port 189 nsew signal output
rlabel metal3 s 0 127032 800 127152 6 o_din0[14]
port 190 nsew signal output
rlabel metal3 s 0 132472 800 132592 6 o_din0[15]
port 191 nsew signal output
rlabel metal2 s 181902 199469 181958 200269 6 o_din0[16]
port 192 nsew signal output
rlabel metal2 s 173806 0 173862 800 6 o_din0[17]
port 193 nsew signal output
rlabel metal2 s 175002 0 175058 800 6 o_din0[18]
port 194 nsew signal output
rlabel metal3 s 197325 138320 198125 138440 6 o_din0[19]
port 195 nsew signal output
rlabel metal3 s 0 24216 800 24336 6 o_din0[1]
port 196 nsew signal output
rlabel metal2 s 179970 0 180026 800 6 o_din0[20]
port 197 nsew signal output
rlabel metal3 s 197325 150152 198125 150272 6 o_din0[21]
port 198 nsew signal output
rlabel metal3 s 197325 156000 198125 156120 6 o_din0[22]
port 199 nsew signal output
rlabel metal2 s 183742 0 183798 800 6 o_din0[23]
port 200 nsew signal output
rlabel metal2 s 189722 199469 189778 200269 6 o_din0[24]
port 201 nsew signal output
rlabel metal2 s 187514 0 187570 800 6 o_din0[25]
port 202 nsew signal output
rlabel metal2 s 188710 0 188766 800 6 o_din0[26]
port 203 nsew signal output
rlabel metal3 s 0 186600 800 186720 6 o_din0[27]
port 204 nsew signal output
rlabel metal2 s 193586 199469 193642 200269 6 o_din0[28]
port 205 nsew signal output
rlabel metal3 s 197325 179528 198125 179648 6 o_din0[29]
port 206 nsew signal output
rlabel metal3 s 0 34960 800 35080 6 o_din0[2]
port 207 nsew signal output
rlabel metal2 s 197450 199469 197506 200269 6 o_din0[30]
port 208 nsew signal output
rlabel metal2 s 197450 0 197506 800 6 o_din0[31]
port 209 nsew signal output
rlabel metal2 s 146390 0 146446 800 6 o_din0[3]
port 210 nsew signal output
rlabel metal2 s 162490 199469 162546 200269 6 o_din0[4]
port 211 nsew signal output
rlabel metal2 s 151358 0 151414 800 6 o_din0[5]
port 212 nsew signal output
rlabel metal2 s 155038 0 155094 800 6 o_din0[6]
port 213 nsew signal output
rlabel metal2 s 169022 199469 169078 200269 6 o_din0[7]
port 214 nsew signal output
rlabel metal3 s 0 94528 800 94648 6 o_din0[8]
port 215 nsew signal output
rlabel metal3 s 0 99968 800 100088 6 o_din0[9]
port 216 nsew signal output
rlabel metal2 s 138846 0 138902 800 6 o_din0_1[0]
port 217 nsew signal output
rlabel metal2 s 161294 0 161350 800 6 o_din0_1[10]
port 218 nsew signal output
rlabel metal3 s 0 110848 800 110968 6 o_din0_1[11]
port 219 nsew signal output
rlabel metal2 s 165066 0 165122 800 6 o_din0_1[12]
port 220 nsew signal output
rlabel metal2 s 168746 0 168802 800 6 o_din0_1[13]
port 221 nsew signal output
rlabel metal3 s 197325 97112 198125 97232 6 o_din0_1[14]
port 222 nsew signal output
rlabel metal2 s 172518 0 172574 800 6 o_din0_1[15]
port 223 nsew signal output
rlabel metal2 s 180614 199469 180670 200269 6 o_din0_1[16]
port 224 nsew signal output
rlabel metal3 s 197325 114792 198125 114912 6 o_din0_1[17]
port 225 nsew signal output
rlabel metal2 s 184570 199469 184626 200269 6 o_din0_1[18]
port 226 nsew signal output
rlabel metal3 s 0 137912 800 138032 6 o_din0_1[19]
port 227 nsew signal output
rlabel metal3 s 197325 26392 198125 26512 6 o_din0_1[1]
port 228 nsew signal output
rlabel metal3 s 0 143352 800 143472 6 o_din0_1[20]
port 229 nsew signal output
rlabel metal2 s 181258 0 181314 800 6 o_din0_1[21]
port 230 nsew signal output
rlabel metal2 s 185858 199469 185914 200269 6 o_din0_1[22]
port 231 nsew signal output
rlabel metal2 s 188434 199469 188490 200269 6 o_din0_1[23]
port 232 nsew signal output
rlabel metal2 s 184938 0 184994 800 6 o_din0_1[24]
port 233 nsew signal output
rlabel metal2 s 186226 0 186282 800 6 o_din0_1[25]
port 234 nsew signal output
rlabel metal3 s 197325 167832 198125 167952 6 o_din0_1[26]
port 235 nsew signal output
rlabel metal3 s 197325 173680 198125 173800 6 o_din0_1[27]
port 236 nsew signal output
rlabel metal2 s 193678 0 193734 800 6 o_din0_1[28]
port 237 nsew signal output
rlabel metal2 s 194966 0 195022 800 6 o_din0_1[29]
port 238 nsew signal output
rlabel metal3 s 0 29656 800 29776 6 o_din0_1[2]
port 239 nsew signal output
rlabel metal3 s 0 192040 800 192160 6 o_din0_1[30]
port 240 nsew signal output
rlabel metal3 s 197325 197208 198125 197328 6 o_din0_1[31]
port 241 nsew signal output
rlabel metal3 s 197325 44072 198125 44192 6 o_din0_1[3]
port 242 nsew signal output
rlabel metal3 s 0 56720 800 56840 6 o_din0_1[4]
port 243 nsew signal output
rlabel metal3 s 0 62024 800 62144 6 o_din0_1[5]
port 244 nsew signal output
rlabel metal2 s 153842 0 153898 800 6 o_din0_1[6]
port 245 nsew signal output
rlabel metal2 s 167734 199469 167790 200269 6 o_din0_1[7]
port 246 nsew signal output
rlabel metal3 s 0 89088 800 89208 6 o_din0_1[8]
port 247 nsew signal output
rlabel metal3 s 197325 79432 198125 79552 6 o_din0_1[9]
port 248 nsew signal output
rlabel metal3 s 197325 8712 198125 8832 6 o_waddr0[0]
port 249 nsew signal output
rlabel metal2 s 154762 199469 154818 200269 6 o_waddr0[1]
port 250 nsew signal output
rlabel metal2 s 156050 199469 156106 200269 6 o_waddr0[2]
port 251 nsew signal output
rlabel metal2 s 147586 0 147642 800 6 o_waddr0[3]
port 252 nsew signal output
rlabel metal3 s 197325 55768 198125 55888 6 o_waddr0[4]
port 253 nsew signal output
rlabel metal2 s 166446 199469 166502 200269 6 o_waddr0[5]
port 254 nsew signal output
rlabel metal2 s 156326 0 156382 800 6 o_waddr0[6]
port 255 nsew signal output
rlabel metal3 s 0 83784 800 83904 6 o_waddr0[7]
port 256 nsew signal output
rlabel metal2 s 160098 0 160154 800 6 o_waddr0[8]
port 257 nsew signal output
rlabel metal2 s 150898 199469 150954 200269 6 o_waddr0_1[0]
port 258 nsew signal output
rlabel metal3 s 197325 32240 198125 32360 6 o_waddr0_1[1]
port 259 nsew signal output
rlabel metal3 s 0 40400 800 40520 6 o_waddr0_1[2]
port 260 nsew signal output
rlabel metal2 s 159914 199469 159970 200269 6 o_waddr0_1[3]
port 261 nsew signal output
rlabel metal2 s 163778 199469 163834 200269 6 o_waddr0_1[4]
port 262 nsew signal output
rlabel metal2 s 165066 199469 165122 200269 6 o_waddr0_1[5]
port 263 nsew signal output
rlabel metal3 s 197325 61752 198125 61872 6 o_waddr0_1[6]
port 264 nsew signal output
rlabel metal3 s 0 78344 800 78464 6 o_waddr0_1[7]
port 265 nsew signal output
rlabel metal3 s 197325 67600 198125 67720 6 o_waddr0_1[8]
port 266 nsew signal output
rlabel metal2 s 149610 199469 149666 200269 6 o_web0
port 267 nsew signal output
rlabel metal3 s 0 13336 800 13456 6 o_web0_1
port 268 nsew signal output
rlabel metal3 s 197325 14560 198125 14680 6 o_wmask0[0]
port 269 nsew signal output
rlabel metal2 s 141330 0 141386 800 6 o_wmask0[1]
port 270 nsew signal output
rlabel metal2 s 157338 199469 157394 200269 6 o_wmask0[2]
port 271 nsew signal output
rlabel metal2 s 161202 199469 161258 200269 6 o_wmask0[3]
port 272 nsew signal output
rlabel metal2 s 152186 199469 152242 200269 6 o_wmask0_1[0]
port 273 nsew signal output
rlabel metal2 s 140134 0 140190 800 6 o_wmask0_1[1]
port 274 nsew signal output
rlabel metal2 s 145102 0 145158 800 6 o_wmask0_1[2]
port 275 nsew signal output
rlabel metal3 s 0 45840 800 45960 6 o_wmask0_1[3]
port 276 nsew signal output
rlabel metal3 s 0 18776 800 18896 6 rst_i
port 277 nsew signal input
rlabel metal4 s 4208 2128 4528 198064 6 vccd1
port 278 nsew power input
rlabel metal4 s 34928 2128 35248 198064 6 vccd1
port 278 nsew power input
rlabel metal4 s 65648 2128 65968 198064 6 vccd1
port 278 nsew power input
rlabel metal4 s 96368 2128 96688 198064 6 vccd1
port 278 nsew power input
rlabel metal4 s 127088 2128 127408 198064 6 vccd1
port 278 nsew power input
rlabel metal4 s 157808 2128 158128 198064 6 vccd1
port 278 nsew power input
rlabel metal4 s 188528 2128 188848 198064 6 vccd1
port 278 nsew power input
rlabel metal4 s 19568 2128 19888 198064 6 vssd1
port 279 nsew ground input
rlabel metal4 s 50288 2128 50608 198064 6 vssd1
port 279 nsew ground input
rlabel metal4 s 81008 2128 81328 198064 6 vssd1
port 279 nsew ground input
rlabel metal4 s 111728 2128 112048 198064 6 vssd1
port 279 nsew ground input
rlabel metal4 s 142448 2128 142768 198064 6 vssd1
port 279 nsew ground input
rlabel metal4 s 173168 2128 173488 198064 6 vssd1
port 279 nsew ground input
rlabel metal2 s 570 0 626 800 6 wb_clk_i
port 280 nsew signal input
rlabel metal2 s 1766 0 1822 800 6 wb_rst_i
port 281 nsew signal input
rlabel metal2 s 3054 0 3110 800 6 wbs_ack_o
port 282 nsew signal output
rlabel metal2 s 8022 0 8078 800 6 wbs_adr_i[0]
port 283 nsew signal input
rlabel metal2 s 50342 0 50398 800 6 wbs_adr_i[10]
port 284 nsew signal input
rlabel metal2 s 54114 0 54170 800 6 wbs_adr_i[11]
port 285 nsew signal input
rlabel metal2 s 57886 0 57942 800 6 wbs_adr_i[12]
port 286 nsew signal input
rlabel metal2 s 61566 0 61622 800 6 wbs_adr_i[13]
port 287 nsew signal input
rlabel metal2 s 65338 0 65394 800 6 wbs_adr_i[14]
port 288 nsew signal input
rlabel metal2 s 69110 0 69166 800 6 wbs_adr_i[15]
port 289 nsew signal input
rlabel metal2 s 72790 0 72846 800 6 wbs_adr_i[16]
port 290 nsew signal input
rlabel metal2 s 76562 0 76618 800 6 wbs_adr_i[17]
port 291 nsew signal input
rlabel metal2 s 80334 0 80390 800 6 wbs_adr_i[18]
port 292 nsew signal input
rlabel metal2 s 84014 0 84070 800 6 wbs_adr_i[19]
port 293 nsew signal input
rlabel metal2 s 12990 0 13046 800 6 wbs_adr_i[1]
port 294 nsew signal input
rlabel metal2 s 87786 0 87842 800 6 wbs_adr_i[20]
port 295 nsew signal input
rlabel metal2 s 91466 0 91522 800 6 wbs_adr_i[21]
port 296 nsew signal input
rlabel metal2 s 95238 0 95294 800 6 wbs_adr_i[22]
port 297 nsew signal input
rlabel metal2 s 99010 0 99066 800 6 wbs_adr_i[23]
port 298 nsew signal input
rlabel metal2 s 102690 0 102746 800 6 wbs_adr_i[24]
port 299 nsew signal input
rlabel metal2 s 106462 0 106518 800 6 wbs_adr_i[25]
port 300 nsew signal input
rlabel metal2 s 110234 0 110290 800 6 wbs_adr_i[26]
port 301 nsew signal input
rlabel metal2 s 113914 0 113970 800 6 wbs_adr_i[27]
port 302 nsew signal input
rlabel metal2 s 117686 0 117742 800 6 wbs_adr_i[28]
port 303 nsew signal input
rlabel metal2 s 121458 0 121514 800 6 wbs_adr_i[29]
port 304 nsew signal input
rlabel metal2 s 17958 0 18014 800 6 wbs_adr_i[2]
port 305 nsew signal input
rlabel metal2 s 125138 0 125194 800 6 wbs_adr_i[30]
port 306 nsew signal input
rlabel metal2 s 128910 0 128966 800 6 wbs_adr_i[31]
port 307 nsew signal input
rlabel metal2 s 22926 0 22982 800 6 wbs_adr_i[3]
port 308 nsew signal input
rlabel metal2 s 27986 0 28042 800 6 wbs_adr_i[4]
port 309 nsew signal input
rlabel metal2 s 31666 0 31722 800 6 wbs_adr_i[5]
port 310 nsew signal input
rlabel metal2 s 35438 0 35494 800 6 wbs_adr_i[6]
port 311 nsew signal input
rlabel metal2 s 39118 0 39174 800 6 wbs_adr_i[7]
port 312 nsew signal input
rlabel metal2 s 42890 0 42946 800 6 wbs_adr_i[8]
port 313 nsew signal input
rlabel metal2 s 46662 0 46718 800 6 wbs_adr_i[9]
port 314 nsew signal input
rlabel metal2 s 4250 0 4306 800 6 wbs_cyc_i
port 315 nsew signal input
rlabel metal2 s 9218 0 9274 800 6 wbs_dat_i[0]
port 316 nsew signal input
rlabel metal2 s 51630 0 51686 800 6 wbs_dat_i[10]
port 317 nsew signal input
rlabel metal2 s 55402 0 55458 800 6 wbs_dat_i[11]
port 318 nsew signal input
rlabel metal2 s 59082 0 59138 800 6 wbs_dat_i[12]
port 319 nsew signal input
rlabel metal2 s 62854 0 62910 800 6 wbs_dat_i[13]
port 320 nsew signal input
rlabel metal2 s 66626 0 66682 800 6 wbs_dat_i[14]
port 321 nsew signal input
rlabel metal2 s 70306 0 70362 800 6 wbs_dat_i[15]
port 322 nsew signal input
rlabel metal2 s 74078 0 74134 800 6 wbs_dat_i[16]
port 323 nsew signal input
rlabel metal2 s 77758 0 77814 800 6 wbs_dat_i[17]
port 324 nsew signal input
rlabel metal2 s 81530 0 81586 800 6 wbs_dat_i[18]
port 325 nsew signal input
rlabel metal2 s 85302 0 85358 800 6 wbs_dat_i[19]
port 326 nsew signal input
rlabel metal2 s 14278 0 14334 800 6 wbs_dat_i[1]
port 327 nsew signal input
rlabel metal2 s 88982 0 89038 800 6 wbs_dat_i[20]
port 328 nsew signal input
rlabel metal2 s 92754 0 92810 800 6 wbs_dat_i[21]
port 329 nsew signal input
rlabel metal2 s 96526 0 96582 800 6 wbs_dat_i[22]
port 330 nsew signal input
rlabel metal2 s 100206 0 100262 800 6 wbs_dat_i[23]
port 331 nsew signal input
rlabel metal2 s 103978 0 104034 800 6 wbs_dat_i[24]
port 332 nsew signal input
rlabel metal2 s 107750 0 107806 800 6 wbs_dat_i[25]
port 333 nsew signal input
rlabel metal2 s 111430 0 111486 800 6 wbs_dat_i[26]
port 334 nsew signal input
rlabel metal2 s 115202 0 115258 800 6 wbs_dat_i[27]
port 335 nsew signal input
rlabel metal2 s 118882 0 118938 800 6 wbs_dat_i[28]
port 336 nsew signal input
rlabel metal2 s 122654 0 122710 800 6 wbs_dat_i[29]
port 337 nsew signal input
rlabel metal2 s 19246 0 19302 800 6 wbs_dat_i[2]
port 338 nsew signal input
rlabel metal2 s 126426 0 126482 800 6 wbs_dat_i[30]
port 339 nsew signal input
rlabel metal2 s 130106 0 130162 800 6 wbs_dat_i[31]
port 340 nsew signal input
rlabel metal2 s 24214 0 24270 800 6 wbs_dat_i[3]
port 341 nsew signal input
rlabel metal2 s 29182 0 29238 800 6 wbs_dat_i[4]
port 342 nsew signal input
rlabel metal2 s 32954 0 33010 800 6 wbs_dat_i[5]
port 343 nsew signal input
rlabel metal2 s 36634 0 36690 800 6 wbs_dat_i[6]
port 344 nsew signal input
rlabel metal2 s 40406 0 40462 800 6 wbs_dat_i[7]
port 345 nsew signal input
rlabel metal2 s 44178 0 44234 800 6 wbs_dat_i[8]
port 346 nsew signal input
rlabel metal2 s 47858 0 47914 800 6 wbs_dat_i[9]
port 347 nsew signal input
rlabel metal2 s 10506 0 10562 800 6 wbs_dat_o[0]
port 348 nsew signal output
rlabel metal2 s 52826 0 52882 800 6 wbs_dat_o[10]
port 349 nsew signal output
rlabel metal2 s 56598 0 56654 800 6 wbs_dat_o[11]
port 350 nsew signal output
rlabel metal2 s 60370 0 60426 800 6 wbs_dat_o[12]
port 351 nsew signal output
rlabel metal2 s 64050 0 64106 800 6 wbs_dat_o[13]
port 352 nsew signal output
rlabel metal2 s 67822 0 67878 800 6 wbs_dat_o[14]
port 353 nsew signal output
rlabel metal2 s 71594 0 71650 800 6 wbs_dat_o[15]
port 354 nsew signal output
rlabel metal2 s 75274 0 75330 800 6 wbs_dat_o[16]
port 355 nsew signal output
rlabel metal2 s 79046 0 79102 800 6 wbs_dat_o[17]
port 356 nsew signal output
rlabel metal2 s 82818 0 82874 800 6 wbs_dat_o[18]
port 357 nsew signal output
rlabel metal2 s 86498 0 86554 800 6 wbs_dat_o[19]
port 358 nsew signal output
rlabel metal2 s 15474 0 15530 800 6 wbs_dat_o[1]
port 359 nsew signal output
rlabel metal2 s 90270 0 90326 800 6 wbs_dat_o[20]
port 360 nsew signal output
rlabel metal2 s 94042 0 94098 800 6 wbs_dat_o[21]
port 361 nsew signal output
rlabel metal2 s 97722 0 97778 800 6 wbs_dat_o[22]
port 362 nsew signal output
rlabel metal2 s 101494 0 101550 800 6 wbs_dat_o[23]
port 363 nsew signal output
rlabel metal2 s 105174 0 105230 800 6 wbs_dat_o[24]
port 364 nsew signal output
rlabel metal2 s 108946 0 109002 800 6 wbs_dat_o[25]
port 365 nsew signal output
rlabel metal2 s 112718 0 112774 800 6 wbs_dat_o[26]
port 366 nsew signal output
rlabel metal2 s 116398 0 116454 800 6 wbs_dat_o[27]
port 367 nsew signal output
rlabel metal2 s 120170 0 120226 800 6 wbs_dat_o[28]
port 368 nsew signal output
rlabel metal2 s 123942 0 123998 800 6 wbs_dat_o[29]
port 369 nsew signal output
rlabel metal2 s 20442 0 20498 800 6 wbs_dat_o[2]
port 370 nsew signal output
rlabel metal2 s 127622 0 127678 800 6 wbs_dat_o[30]
port 371 nsew signal output
rlabel metal2 s 131394 0 131450 800 6 wbs_dat_o[31]
port 372 nsew signal output
rlabel metal2 s 25410 0 25466 800 6 wbs_dat_o[3]
port 373 nsew signal output
rlabel metal2 s 30470 0 30526 800 6 wbs_dat_o[4]
port 374 nsew signal output
rlabel metal2 s 34150 0 34206 800 6 wbs_dat_o[5]
port 375 nsew signal output
rlabel metal2 s 37922 0 37978 800 6 wbs_dat_o[6]
port 376 nsew signal output
rlabel metal2 s 41694 0 41750 800 6 wbs_dat_o[7]
port 377 nsew signal output
rlabel metal2 s 45374 0 45430 800 6 wbs_dat_o[8]
port 378 nsew signal output
rlabel metal2 s 49146 0 49202 800 6 wbs_dat_o[9]
port 379 nsew signal output
rlabel metal2 s 11702 0 11758 800 6 wbs_sel_i[0]
port 380 nsew signal input
rlabel metal2 s 16762 0 16818 800 6 wbs_sel_i[1]
port 381 nsew signal input
rlabel metal2 s 21730 0 21786 800 6 wbs_sel_i[2]
port 382 nsew signal input
rlabel metal2 s 26698 0 26754 800 6 wbs_sel_i[3]
port 383 nsew signal input
rlabel metal2 s 5538 0 5594 800 6 wbs_stb_i
port 384 nsew signal input
rlabel metal2 s 6734 0 6790 800 6 wbs_we_i
port 385 nsew signal input
<< properties >>
string LEFclass BLOCK
string FIXED_BBOX 0 0 198125 200269
string LEFview TRUE
string GDS_FILE /local/home/roman/projects/opencircuitdesign/shuttle5/caravel_mpw/openlane/user_proj/runs/user_proj/results/magic/user_proj.gds
string GDS_END 97554168
string GDS_START 1460416
<< end >>

