VERSION 5.7 ;
  NOWIREEXTENSIONATPIN ON ;
  DIVIDERCHAR "/" ;
  BUSBITCHARS "[]" ;
MACRO user_proj
  CLASS BLOCK ;
  FOREIGN user_proj ;
  ORIGIN 0.000 0.000 ;
  SIZE 997.120 BY 1007.840 ;
  PIN clk_i
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 779.330 0.000 779.610 4.000 ;
    END
  END clk_i
  PIN i_dout0[0]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 793.590 0.000 793.870 4.000 ;
    END
  END i_dout0[0]
  PIN i_dout0[10]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 514.800 4.000 515.400 ;
    END
  END i_dout0[10]
  PIN i_dout0[11]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 830.390 1003.840 830.670 1007.840 ;
    END
  END i_dout0[11]
  PIN i_dout0[12]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 836.830 1003.840 837.110 1007.840 ;
    END
  END i_dout0[12]
  PIN i_dout0[13]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 580.080 4.000 580.680 ;
    END
  END i_dout0[13]
  PIN i_dout0[14]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 993.120 490.320 997.120 490.920 ;
    END
  END i_dout0[14]
  PIN i_dout0[15]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 993.120 569.880 997.120 570.480 ;
    END
  END i_dout0[15]
  PIN i_dout0[16]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 624.280 4.000 624.880 ;
    END
  END i_dout0[16]
  PIN i_dout0[17]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 993.120 622.920 997.120 623.520 ;
    END
  END i_dout0[17]
  PIN i_dout0[18]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 667.800 4.000 668.400 ;
    END
  END i_dout0[18]
  PIN i_dout0[19]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 893.410 1003.840 893.690 1007.840 ;
    END
  END i_dout0[19]
  PIN i_dout0[1]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 76.200 4.000 76.800 ;
    END
  END i_dout0[1]
  PIN i_dout0[20]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 905.830 1003.840 906.110 1007.840 ;
    END
  END i_dout0[20]
  PIN i_dout0[21]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 936.190 0.000 936.470 4.000 ;
    END
  END i_dout0[21]
  PIN i_dout0[22]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 799.040 4.000 799.640 ;
    END
  END i_dout0[22]
  PIN i_dout0[23]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 931.130 1003.840 931.410 1007.840 ;
    END
  END i_dout0[23]
  PIN i_dout0[24]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 993.120 861.600 997.120 862.200 ;
    END
  END i_dout0[24]
  PIN i_dout0[25]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 943.550 1003.840 943.830 1007.840 ;
    END
  END i_dout0[25]
  PIN i_dout0[26]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 865.000 4.000 865.600 ;
    END
  END i_dout0[26]
  PIN i_dout0[27]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 886.760 4.000 887.360 ;
    END
  END i_dout0[27]
  PIN i_dout0[28]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 993.120 941.160 997.120 941.760 ;
    END
  END i_dout0[28]
  PIN i_dout0[29]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 993.230 0.000 993.510 4.000 ;
    END
  END i_dout0[29]
  PIN i_dout0[2]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 993.120 172.080 997.120 172.680 ;
    END
  END i_dout0[2]
  PIN i_dout0[30]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 974.480 4.000 975.080 ;
    END
  END i_dout0[30]
  PIN i_dout0[31]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 993.120 994.200 997.120 994.800 ;
    END
  END i_dout0[31]
  PIN i_dout0[3]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 993.120 251.640 997.120 252.240 ;
    END
  END i_dout0[3]
  PIN i_dout0[4]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 993.120 331.200 997.120 331.800 ;
    END
  END i_dout0[4]
  PIN i_dout0[5]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 774.270 1003.840 774.550 1007.840 ;
    END
  END i_dout0[5]
  PIN i_dout0[6]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 361.120 4.000 361.720 ;
    END
  END i_dout0[6]
  PIN i_dout0[7]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 850.630 0.000 850.910 4.000 ;
    END
  END i_dout0[7]
  PIN i_dout0[8]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 805.550 1003.840 805.830 1007.840 ;
    END
  END i_dout0[8]
  PIN i_dout0[9]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 893.410 0.000 893.690 4.000 ;
    END
  END i_dout0[9]
  PIN i_dout0_1[0]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 800.950 0.000 801.230 4.000 ;
    END
  END i_dout0_1[0]
  PIN i_dout0_1[10]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 993.120 437.280 997.120 437.880 ;
    END
  END i_dout0_1[10]
  PIN i_dout0_1[11]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 536.560 4.000 537.160 ;
    END
  END i_dout0_1[11]
  PIN i_dout0_1[12]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 915.030 0.000 915.310 4.000 ;
    END
  END i_dout0_1[12]
  PIN i_dout0_1[13]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 843.270 1003.840 843.550 1007.840 ;
    END
  END i_dout0_1[13]
  PIN i_dout0_1[14]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 929.290 0.000 929.570 4.000 ;
    END
  END i_dout0_1[14]
  PIN i_dout0_1[15]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 993.120 543.360 997.120 543.960 ;
    END
  END i_dout0_1[15]
  PIN i_dout0_1[16]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 601.840 4.000 602.440 ;
    END
  END i_dout0_1[16]
  PIN i_dout0_1[17]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 646.040 4.000 646.640 ;
    END
  END i_dout0_1[17]
  PIN i_dout0_1[18]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 886.970 1003.840 887.250 1007.840 ;
    END
  END i_dout0_1[18]
  PIN i_dout0_1[19]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 993.120 675.960 997.120 676.560 ;
    END
  END i_dout0_1[19]
  PIN i_dout0_1[1]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 807.850 0.000 808.130 4.000 ;
    END
  END i_dout0_1[1]
  PIN i_dout0_1[20]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 993.120 702.480 997.120 703.080 ;
    END
  END i_dout0_1[20]
  PIN i_dout0_1[21]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 777.280 4.000 777.880 ;
    END
  END i_dout0_1[21]
  PIN i_dout0_1[22]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 918.250 1003.840 918.530 1007.840 ;
    END
  END i_dout0_1[22]
  PIN i_dout0_1[23]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 993.120 782.040 997.120 782.640 ;
    END
  END i_dout0_1[23]
  PIN i_dout0_1[24]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 993.120 835.080 997.120 835.680 ;
    END
  END i_dout0_1[24]
  PIN i_dout0_1[25]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 950.450 0.000 950.730 4.000 ;
    END
  END i_dout0_1[25]
  PIN i_dout0_1[26]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 957.810 0.000 958.090 4.000 ;
    END
  END i_dout0_1[26]
  PIN i_dout0_1[27]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 993.120 914.640 997.120 915.240 ;
    END
  END i_dout0_1[27]
  PIN i_dout0_1[28]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 978.970 0.000 979.250 4.000 ;
    END
  END i_dout0_1[28]
  PIN i_dout0_1[29]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 930.960 4.000 931.560 ;
    END
  END i_dout0_1[29]
  PIN i_dout0_1[2]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 815.210 0.000 815.490 4.000 ;
    END
  END i_dout0_1[2]
  PIN i_dout0_1[30]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 952.720 4.000 953.320 ;
    END
  END i_dout0_1[30]
  PIN i_dout0_1[31]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 987.250 1003.840 987.530 1007.840 ;
    END
  END i_dout0_1[31]
  PIN i_dout0_1[3]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 829.470 0.000 829.750 4.000 ;
    END
  END i_dout0_1[3]
  PIN i_dout0_1[4]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 755.410 1003.840 755.690 1007.840 ;
    END
  END i_dout0_1[4]
  PIN i_dout0_1[5]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 273.400 4.000 274.000 ;
    END
  END i_dout0_1[5]
  PIN i_dout0_1[6]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 339.360 4.000 339.960 ;
    END
  END i_dout0_1[6]
  PIN i_dout0_1[7]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 799.110 1003.840 799.390 1007.840 ;
    END
  END i_dout0_1[7]
  PIN i_dout0_1[8]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 448.840 4.000 449.440 ;
    END
  END i_dout0_1[8]
  PIN i_dout0_1[9]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 886.510 0.000 886.790 4.000 ;
    END
  END i_dout0_1[9]
  PIN io_in[0]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 2.850 1003.840 3.130 1007.840 ;
    END
  END io_in[0]
  PIN io_in[10]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 190.990 1003.840 191.270 1007.840 ;
    END
  END io_in[10]
  PIN io_in[11]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 209.390 1003.840 209.670 1007.840 ;
    END
  END io_in[11]
  PIN io_in[12]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 228.250 1003.840 228.530 1007.840 ;
    END
  END io_in[12]
  PIN io_in[13]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 247.110 1003.840 247.390 1007.840 ;
    END
  END io_in[13]
  PIN io_in[14]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 265.970 1003.840 266.250 1007.840 ;
    END
  END io_in[14]
  PIN io_in[15]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 284.830 1003.840 285.110 1007.840 ;
    END
  END io_in[15]
  PIN io_in[16]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 303.690 1003.840 303.970 1007.840 ;
    END
  END io_in[16]
  PIN io_in[17]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 322.550 1003.840 322.830 1007.840 ;
    END
  END io_in[17]
  PIN io_in[18]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 341.410 1003.840 341.690 1007.840 ;
    END
  END io_in[18]
  PIN io_in[19]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 360.270 1003.840 360.550 1007.840 ;
    END
  END io_in[19]
  PIN io_in[1]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 21.250 1003.840 21.530 1007.840 ;
    END
  END io_in[1]
  PIN io_in[20]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 379.130 1003.840 379.410 1007.840 ;
    END
  END io_in[20]
  PIN io_in[21]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 397.990 1003.840 398.270 1007.840 ;
    END
  END io_in[21]
  PIN io_in[22]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 416.390 1003.840 416.670 1007.840 ;
    END
  END io_in[22]
  PIN io_in[23]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 435.250 1003.840 435.530 1007.840 ;
    END
  END io_in[23]
  PIN io_in[24]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 454.110 1003.840 454.390 1007.840 ;
    END
  END io_in[24]
  PIN io_in[25]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 472.970 1003.840 473.250 1007.840 ;
    END
  END io_in[25]
  PIN io_in[26]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 491.830 1003.840 492.110 1007.840 ;
    END
  END io_in[26]
  PIN io_in[27]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 510.690 1003.840 510.970 1007.840 ;
    END
  END io_in[27]
  PIN io_in[28]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 529.550 1003.840 529.830 1007.840 ;
    END
  END io_in[28]
  PIN io_in[29]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 548.410 1003.840 548.690 1007.840 ;
    END
  END io_in[29]
  PIN io_in[2]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 40.110 1003.840 40.390 1007.840 ;
    END
  END io_in[2]
  PIN io_in[30]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 567.270 1003.840 567.550 1007.840 ;
    END
  END io_in[30]
  PIN io_in[31]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 586.130 1003.840 586.410 1007.840 ;
    END
  END io_in[31]
  PIN io_in[32]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 604.530 1003.840 604.810 1007.840 ;
    END
  END io_in[32]
  PIN io_in[33]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 623.390 1003.840 623.670 1007.840 ;
    END
  END io_in[33]
  PIN io_in[34]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 642.250 1003.840 642.530 1007.840 ;
    END
  END io_in[34]
  PIN io_in[35]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 661.110 1003.840 661.390 1007.840 ;
    END
  END io_in[35]
  PIN io_in[36]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 679.970 1003.840 680.250 1007.840 ;
    END
  END io_in[36]
  PIN io_in[37]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 698.830 1003.840 699.110 1007.840 ;
    END
  END io_in[37]
  PIN io_in[3]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 58.970 1003.840 59.250 1007.840 ;
    END
  END io_in[3]
  PIN io_in[4]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 77.830 1003.840 78.110 1007.840 ;
    END
  END io_in[4]
  PIN io_in[5]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 96.690 1003.840 96.970 1007.840 ;
    END
  END io_in[5]
  PIN io_in[6]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 115.550 1003.840 115.830 1007.840 ;
    END
  END io_in[6]
  PIN io_in[7]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 134.410 1003.840 134.690 1007.840 ;
    END
  END io_in[7]
  PIN io_in[8]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 153.270 1003.840 153.550 1007.840 ;
    END
  END io_in[8]
  PIN io_in[9]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 172.130 1003.840 172.410 1007.840 ;
    END
  END io_in[9]
  PIN io_oeb[0]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 8.830 1003.840 9.110 1007.840 ;
    END
  END io_oeb[0]
  PIN io_oeb[10]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 196.970 1003.840 197.250 1007.840 ;
    END
  END io_oeb[10]
  PIN io_oeb[11]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 215.830 1003.840 216.110 1007.840 ;
    END
  END io_oeb[11]
  PIN io_oeb[12]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 234.690 1003.840 234.970 1007.840 ;
    END
  END io_oeb[12]
  PIN io_oeb[13]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 253.550 1003.840 253.830 1007.840 ;
    END
  END io_oeb[13]
  PIN io_oeb[14]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 272.410 1003.840 272.690 1007.840 ;
    END
  END io_oeb[14]
  PIN io_oeb[15]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 291.270 1003.840 291.550 1007.840 ;
    END
  END io_oeb[15]
  PIN io_oeb[16]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 310.130 1003.840 310.410 1007.840 ;
    END
  END io_oeb[16]
  PIN io_oeb[17]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 328.990 1003.840 329.270 1007.840 ;
    END
  END io_oeb[17]
  PIN io_oeb[18]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 347.390 1003.840 347.670 1007.840 ;
    END
  END io_oeb[18]
  PIN io_oeb[19]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 366.250 1003.840 366.530 1007.840 ;
    END
  END io_oeb[19]
  PIN io_oeb[1]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 27.690 1003.840 27.970 1007.840 ;
    END
  END io_oeb[1]
  PIN io_oeb[20]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 385.110 1003.840 385.390 1007.840 ;
    END
  END io_oeb[20]
  PIN io_oeb[21]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 403.970 1003.840 404.250 1007.840 ;
    END
  END io_oeb[21]
  PIN io_oeb[22]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 422.830 1003.840 423.110 1007.840 ;
    END
  END io_oeb[22]
  PIN io_oeb[23]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 441.690 1003.840 441.970 1007.840 ;
    END
  END io_oeb[23]
  PIN io_oeb[24]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 460.550 1003.840 460.830 1007.840 ;
    END
  END io_oeb[24]
  PIN io_oeb[25]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 479.410 1003.840 479.690 1007.840 ;
    END
  END io_oeb[25]
  PIN io_oeb[26]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 498.270 1003.840 498.550 1007.840 ;
    END
  END io_oeb[26]
  PIN io_oeb[27]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 517.130 1003.840 517.410 1007.840 ;
    END
  END io_oeb[27]
  PIN io_oeb[28]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 535.530 1003.840 535.810 1007.840 ;
    END
  END io_oeb[28]
  PIN io_oeb[29]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 554.390 1003.840 554.670 1007.840 ;
    END
  END io_oeb[29]
  PIN io_oeb[2]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 46.550 1003.840 46.830 1007.840 ;
    END
  END io_oeb[2]
  PIN io_oeb[30]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 573.250 1003.840 573.530 1007.840 ;
    END
  END io_oeb[30]
  PIN io_oeb[31]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 592.110 1003.840 592.390 1007.840 ;
    END
  END io_oeb[31]
  PIN io_oeb[32]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 610.970 1003.840 611.250 1007.840 ;
    END
  END io_oeb[32]
  PIN io_oeb[33]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 629.830 1003.840 630.110 1007.840 ;
    END
  END io_oeb[33]
  PIN io_oeb[34]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 648.690 1003.840 648.970 1007.840 ;
    END
  END io_oeb[34]
  PIN io_oeb[35]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 667.550 1003.840 667.830 1007.840 ;
    END
  END io_oeb[35]
  PIN io_oeb[36]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 686.410 1003.840 686.690 1007.840 ;
    END
  END io_oeb[36]
  PIN io_oeb[37]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 705.270 1003.840 705.550 1007.840 ;
    END
  END io_oeb[37]
  PIN io_oeb[3]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 65.410 1003.840 65.690 1007.840 ;
    END
  END io_oeb[3]
  PIN io_oeb[4]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 84.270 1003.840 84.550 1007.840 ;
    END
  END io_oeb[4]
  PIN io_oeb[5]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 103.130 1003.840 103.410 1007.840 ;
    END
  END io_oeb[5]
  PIN io_oeb[6]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 121.990 1003.840 122.270 1007.840 ;
    END
  END io_oeb[6]
  PIN io_oeb[7]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 140.390 1003.840 140.670 1007.840 ;
    END
  END io_oeb[7]
  PIN io_oeb[8]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 159.250 1003.840 159.530 1007.840 ;
    END
  END io_oeb[8]
  PIN io_oeb[9]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 178.110 1003.840 178.390 1007.840 ;
    END
  END io_oeb[9]
  PIN io_out[0]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 15.270 1003.840 15.550 1007.840 ;
    END
  END io_out[0]
  PIN io_out[10]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 203.410 1003.840 203.690 1007.840 ;
    END
  END io_out[10]
  PIN io_out[11]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 222.270 1003.840 222.550 1007.840 ;
    END
  END io_out[11]
  PIN io_out[12]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 241.130 1003.840 241.410 1007.840 ;
    END
  END io_out[12]
  PIN io_out[13]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 259.990 1003.840 260.270 1007.840 ;
    END
  END io_out[13]
  PIN io_out[14]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 278.390 1003.840 278.670 1007.840 ;
    END
  END io_out[14]
  PIN io_out[15]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 297.250 1003.840 297.530 1007.840 ;
    END
  END io_out[15]
  PIN io_out[16]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 316.110 1003.840 316.390 1007.840 ;
    END
  END io_out[16]
  PIN io_out[17]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 334.970 1003.840 335.250 1007.840 ;
    END
  END io_out[17]
  PIN io_out[18]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 353.830 1003.840 354.110 1007.840 ;
    END
  END io_out[18]
  PIN io_out[19]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 372.690 1003.840 372.970 1007.840 ;
    END
  END io_out[19]
  PIN io_out[1]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 34.130 1003.840 34.410 1007.840 ;
    END
  END io_out[1]
  PIN io_out[20]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 391.550 1003.840 391.830 1007.840 ;
    END
  END io_out[20]
  PIN io_out[21]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 410.410 1003.840 410.690 1007.840 ;
    END
  END io_out[21]
  PIN io_out[22]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 429.270 1003.840 429.550 1007.840 ;
    END
  END io_out[22]
  PIN io_out[23]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 448.130 1003.840 448.410 1007.840 ;
    END
  END io_out[23]
  PIN io_out[24]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 466.990 1003.840 467.270 1007.840 ;
    END
  END io_out[24]
  PIN io_out[25]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 485.390 1003.840 485.670 1007.840 ;
    END
  END io_out[25]
  PIN io_out[26]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 504.250 1003.840 504.530 1007.840 ;
    END
  END io_out[26]
  PIN io_out[27]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 523.110 1003.840 523.390 1007.840 ;
    END
  END io_out[27]
  PIN io_out[28]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 541.970 1003.840 542.250 1007.840 ;
    END
  END io_out[28]
  PIN io_out[29]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 560.830 1003.840 561.110 1007.840 ;
    END
  END io_out[29]
  PIN io_out[2]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 52.990 1003.840 53.270 1007.840 ;
    END
  END io_out[2]
  PIN io_out[30]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 579.690 1003.840 579.970 1007.840 ;
    END
  END io_out[30]
  PIN io_out[31]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 598.550 1003.840 598.830 1007.840 ;
    END
  END io_out[31]
  PIN io_out[32]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 617.410 1003.840 617.690 1007.840 ;
    END
  END io_out[32]
  PIN io_out[33]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 636.270 1003.840 636.550 1007.840 ;
    END
  END io_out[33]
  PIN io_out[34]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 655.130 1003.840 655.410 1007.840 ;
    END
  END io_out[34]
  PIN io_out[35]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 673.530 1003.840 673.810 1007.840 ;
    END
  END io_out[35]
  PIN io_out[36]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 692.390 1003.840 692.670 1007.840 ;
    END
  END io_out[36]
  PIN io_out[37]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 711.250 1003.840 711.530 1007.840 ;
    END
  END io_out[37]
  PIN io_out[3]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 71.390 1003.840 71.670 1007.840 ;
    END
  END io_out[3]
  PIN io_out[4]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 90.250 1003.840 90.530 1007.840 ;
    END
  END io_out[4]
  PIN io_out[5]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 109.110 1003.840 109.390 1007.840 ;
    END
  END io_out[5]
  PIN io_out[6]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 127.970 1003.840 128.250 1007.840 ;
    END
  END io_out[6]
  PIN io_out[7]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 146.830 1003.840 147.110 1007.840 ;
    END
  END io_out[7]
  PIN io_out[8]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 165.690 1003.840 165.970 1007.840 ;
    END
  END io_out[8]
  PIN io_out[9]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 184.550 1003.840 184.830 1007.840 ;
    END
  END io_out[9]
  PIN irq[0]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 758.170 0.000 758.450 4.000 ;
    END
  END irq[0]
  PIN irq[1]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 765.070 0.000 765.350 4.000 ;
    END
  END irq[1]
  PIN irq[2]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 772.430 0.000 772.710 4.000 ;
    END
  END irq[2]
  PIN o_csb0
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 10.920 4.000 11.520 ;
    END
  END o_csb0
  PIN o_csb0_1
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 32.680 4.000 33.280 ;
    END
  END o_csb0_1
  PIN o_din0[0]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 993.120 12.960 997.120 13.560 ;
    END
  END o_din0[0]
  PIN o_din0[10]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 824.410 1003.840 824.690 1007.840 ;
    END
  END o_din0[10]
  PIN o_din0[11]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 907.670 0.000 907.950 4.000 ;
    END
  END o_din0[11]
  PIN o_din0[12]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 993.120 463.800 997.120 464.400 ;
    END
  END o_din0[12]
  PIN o_din0[13]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 921.930 0.000 922.210 4.000 ;
    END
  END o_din0[13]
  PIN o_din0[14]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 993.120 516.840 997.120 517.440 ;
    END
  END o_din0[14]
  PIN o_din0[15]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 868.110 1003.840 868.390 1007.840 ;
    END
  END o_din0[15]
  PIN o_din0[16]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 993.120 596.400 997.120 597.000 ;
    END
  END o_din0[16]
  PIN o_din0[17]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 993.120 649.440 997.120 650.040 ;
    END
  END o_din0[17]
  PIN o_din0[18]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 711.320 4.000 711.920 ;
    END
  END o_din0[18]
  PIN o_din0[19]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 899.390 1003.840 899.670 1007.840 ;
    END
  END o_din0[19]
  PIN o_din0[1]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 993.120 92.520 997.120 93.120 ;
    END
  END o_din0[1]
  PIN o_din0[20]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 912.270 1003.840 912.550 1007.840 ;
    END
  END o_din0[20]
  PIN o_din0[21]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 993.120 755.520 997.120 756.120 ;
    END
  END o_din0[21]
  PIN o_din0[22]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 821.480 4.000 822.080 ;
    END
  END o_din0[22]
  PIN o_din0[23]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 937.110 1003.840 937.390 1007.840 ;
    END
  END o_din0[23]
  PIN o_din0[24]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 943.550 0.000 943.830 4.000 ;
    END
  END o_din0[24]
  PIN o_din0[25]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 843.240 4.000 843.840 ;
    END
  END o_din0[25]
  PIN o_din0[26]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 955.970 1003.840 956.250 1007.840 ;
    END
  END o_din0[26]
  PIN o_din0[27]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 962.410 1003.840 962.690 1007.840 ;
    END
  END o_din0[27]
  PIN o_din0[28]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 986.330 0.000 986.610 4.000 ;
    END
  END o_din0[28]
  PIN o_din0[29]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 974.830 1003.840 975.110 1007.840 ;
    END
  END o_din0[29]
  PIN o_din0[2]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 163.920 4.000 164.520 ;
    END
  END o_din0[2]
  PIN o_din0[30]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 981.270 1003.840 981.550 1007.840 ;
    END
  END o_din0[30]
  PIN o_din0[31]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 996.240 4.000 996.840 ;
    END
  END o_din0[31]
  PIN o_din0[3]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 207.440 4.000 208.040 ;
    END
  END o_din0[3]
  PIN o_din0[4]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 993.120 357.720 997.120 358.320 ;
    END
  END o_din0[4]
  PIN o_din0[5]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 317.600 4.000 318.200 ;
    END
  END o_din0[5]
  PIN o_din0[6]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 404.640 4.000 405.240 ;
    END
  END o_din0[6]
  PIN o_din0[7]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 427.080 4.000 427.680 ;
    END
  END o_din0[7]
  PIN o_din0[8]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 872.250 0.000 872.530 4.000 ;
    END
  END o_din0[8]
  PIN o_din0[9]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 993.120 410.760 997.120 411.360 ;
    END
  END o_din0[9]
  PIN o_din0_1[0]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 730.110 1003.840 730.390 1007.840 ;
    END
  END o_din0_1[0]
  PIN o_din0_1[10]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 817.970 1003.840 818.250 1007.840 ;
    END
  END o_din0_1[10]
  PIN o_din0_1[11]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 900.770 0.000 901.050 4.000 ;
    END
  END o_din0_1[11]
  PIN o_din0_1[12]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 558.320 4.000 558.920 ;
    END
  END o_din0_1[12]
  PIN o_din0_1[13]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 849.250 1003.840 849.530 1007.840 ;
    END
  END o_din0_1[13]
  PIN o_din0_1[14]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 855.690 1003.840 855.970 1007.840 ;
    END
  END o_din0_1[14]
  PIN o_din0_1[15]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 862.130 1003.840 862.410 1007.840 ;
    END
  END o_din0_1[15]
  PIN o_din0_1[16]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 874.550 1003.840 874.830 1007.840 ;
    END
  END o_din0_1[16]
  PIN o_din0_1[17]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 880.530 1003.840 880.810 1007.840 ;
    END
  END o_din0_1[17]
  PIN o_din0_1[18]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 689.560 4.000 690.160 ;
    END
  END o_din0_1[18]
  PIN o_din0_1[19]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 733.760 4.000 734.360 ;
    END
  END o_din0_1[19]
  PIN o_din0_1[1]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 742.530 1003.840 742.810 1007.840 ;
    END
  END o_din0_1[1]
  PIN o_din0_1[20]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 755.520 4.000 756.120 ;
    END
  END o_din0_1[20]
  PIN o_din0_1[21]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 993.120 729.000 997.120 729.600 ;
    END
  END o_din0_1[21]
  PIN o_din0_1[22]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 924.690 1003.840 924.970 1007.840 ;
    END
  END o_din0_1[22]
  PIN o_din0_1[23]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 993.120 808.560 997.120 809.160 ;
    END
  END o_din0_1[23]
  PIN o_din0_1[24]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 993.120 888.120 997.120 888.720 ;
    END
  END o_din0_1[24]
  PIN o_din0_1[25]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 949.530 1003.840 949.810 1007.840 ;
    END
  END o_din0_1[25]
  PIN o_din0_1[26]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 964.710 0.000 964.990 4.000 ;
    END
  END o_din0_1[26]
  PIN o_din0_1[27]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 972.070 0.000 972.350 4.000 ;
    END
  END o_din0_1[27]
  PIN o_din0_1[28]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 908.520 4.000 909.120 ;
    END
  END o_din0_1[28]
  PIN o_din0_1[29]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 968.390 1003.840 968.670 1007.840 ;
    END
  END o_din0_1[29]
  PIN o_din0_1[2]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 142.160 4.000 142.760 ;
    END
  END o_din0_1[2]
  PIN o_din0_1[30]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 993.120 967.680 997.120 968.280 ;
    END
  END o_din0_1[30]
  PIN o_din0_1[31]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 993.690 1003.840 993.970 1007.840 ;
    END
  END o_din0_1[31]
  PIN o_din0_1[3]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 836.370 0.000 836.650 4.000 ;
    END
  END o_din0_1[3]
  PIN o_din0_1[4]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 251.640 4.000 252.240 ;
    END
  END o_din0_1[4]
  PIN o_din0_1[5]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 295.160 4.000 295.760 ;
    END
  END o_din0_1[5]
  PIN o_din0_1[6]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 382.880 4.000 383.480 ;
    END
  END o_din0_1[6]
  PIN o_din0_1[7]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 857.990 0.000 858.270 4.000 ;
    END
  END o_din0_1[7]
  PIN o_din0_1[8]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 811.530 1003.840 811.810 1007.840 ;
    END
  END o_din0_1[8]
  PIN o_din0_1[9]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 492.360 4.000 492.960 ;
    END
  END o_din0_1[9]
  PIN o_waddr0[0]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 993.120 39.480 997.120 40.080 ;
    END
  END o_waddr0[0]
  PIN o_waddr0[1]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 993.120 145.560 997.120 146.160 ;
    END
  END o_waddr0[1]
  PIN o_waddr0[2]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 993.120 225.120 997.120 225.720 ;
    END
  END o_waddr0[2]
  PIN o_waddr0[3]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 748.970 1003.840 749.250 1007.840 ;
    END
  END o_waddr0[3]
  PIN o_waddr0[4]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 767.830 1003.840 768.110 1007.840 ;
    END
  END o_waddr0[4]
  PIN o_waddr0[5]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 780.250 1003.840 780.530 1007.840 ;
    END
  END o_waddr0[5]
  PIN o_waddr0[6]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 793.130 1003.840 793.410 1007.840 ;
    END
  END o_waddr0[6]
  PIN o_waddr0[7]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 864.890 0.000 865.170 4.000 ;
    END
  END o_waddr0[7]
  PIN o_waddr0[8]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 879.150 0.000 879.430 4.000 ;
    END
  END o_waddr0[8]
  PIN o_waddr0_1[0]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 54.440 4.000 55.040 ;
    END
  END o_waddr0_1[0]
  PIN o_waddr0_1[1]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 993.120 119.040 997.120 119.640 ;
    END
  END o_waddr0_1[1]
  PIN o_waddr0_1[2]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 993.120 198.600 997.120 199.200 ;
    END
  END o_waddr0_1[2]
  PIN o_waddr0_1[3]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 993.120 278.160 997.120 278.760 ;
    END
  END o_waddr0_1[3]
  PIN o_waddr0_1[4]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 761.390 1003.840 761.670 1007.840 ;
    END
  END o_waddr0_1[4]
  PIN o_waddr0_1[5]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 843.730 0.000 844.010 4.000 ;
    END
  END o_waddr0_1[5]
  PIN o_waddr0_1[6]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 786.690 1003.840 786.970 1007.840 ;
    END
  END o_waddr0_1[6]
  PIN o_waddr0_1[7]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 993.120 384.240 997.120 384.840 ;
    END
  END o_waddr0_1[7]
  PIN o_waddr0_1[8]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 470.600 4.000 471.200 ;
    END
  END o_waddr0_1[8]
  PIN o_web0
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 786.690 0.000 786.970 4.000 ;
    END
  END o_web0
  PIN o_web0_1
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 717.690 1003.840 717.970 1007.840 ;
    END
  END o_web0_1
  PIN o_wmask0[0]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 736.550 1003.840 736.830 1007.840 ;
    END
  END o_wmask0[0]
  PIN o_wmask0[1]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 120.400 4.000 121.000 ;
    END
  END o_wmask0[1]
  PIN o_wmask0[2]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 822.110 0.000 822.390 4.000 ;
    END
  END o_wmask0[2]
  PIN o_wmask0[3]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 993.120 304.680 997.120 305.280 ;
    END
  END o_wmask0[3]
  PIN o_wmask0_1[0]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 993.120 66.000 997.120 66.600 ;
    END
  END o_wmask0_1[0]
  PIN o_wmask0_1[1]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 97.960 4.000 98.560 ;
    END
  END o_wmask0_1[1]
  PIN o_wmask0_1[2]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 185.680 4.000 186.280 ;
    END
  END o_wmask0_1[2]
  PIN o_wmask0_1[3]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 229.880 4.000 230.480 ;
    END
  END o_wmask0_1[3]
  PIN rst_i
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 724.130 1003.840 724.410 1007.840 ;
    END
  END rst_i
  PIN vccd1
    DIRECTION INPUT ;
    USE POWER ;
    PORT
      LAYER met4 ;
        RECT 21.040 10.640 22.640 995.760 ;
    END
    PORT
      LAYER met4 ;
        RECT 174.640 10.640 176.240 995.760 ;
    END
    PORT
      LAYER met4 ;
        RECT 328.240 10.640 329.840 995.760 ;
    END
    PORT
      LAYER met4 ;
        RECT 481.840 10.640 483.440 995.760 ;
    END
    PORT
      LAYER met4 ;
        RECT 635.440 10.640 637.040 995.760 ;
    END
    PORT
      LAYER met4 ;
        RECT 789.040 10.640 790.640 995.760 ;
    END
    PORT
      LAYER met4 ;
        RECT 942.640 10.640 944.240 995.760 ;
    END
  END vccd1
  PIN vssd1
    DIRECTION INPUT ;
    USE GROUND ;
    PORT
      LAYER met4 ;
        RECT 97.840 10.640 99.440 995.760 ;
    END
    PORT
      LAYER met4 ;
        RECT 251.440 10.640 253.040 995.760 ;
    END
    PORT
      LAYER met4 ;
        RECT 405.040 10.640 406.640 995.760 ;
    END
    PORT
      LAYER met4 ;
        RECT 558.640 10.640 560.240 995.760 ;
    END
    PORT
      LAYER met4 ;
        RECT 712.240 10.640 713.840 995.760 ;
    END
    PORT
      LAYER met4 ;
        RECT 865.840 10.640 867.440 995.760 ;
    END
  END vssd1
  PIN wb_clk_i
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 3.310 0.000 3.590 4.000 ;
    END
  END wb_clk_i
  PIN wb_rst_i
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 10.210 0.000 10.490 4.000 ;
    END
  END wb_rst_i
  PIN wbs_ack_o
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 17.110 0.000 17.390 4.000 ;
    END
  END wbs_ack_o
  PIN wbs_adr_i[0]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 45.630 0.000 45.910 4.000 ;
    END
  END wbs_adr_i[0]
  PIN wbs_adr_i[10]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 288.050 0.000 288.330 4.000 ;
    END
  END wbs_adr_i[10]
  PIN wbs_adr_i[11]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 309.210 0.000 309.490 4.000 ;
    END
  END wbs_adr_i[11]
  PIN wbs_adr_i[12]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 330.830 0.000 331.110 4.000 ;
    END
  END wbs_adr_i[12]
  PIN wbs_adr_i[13]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 351.990 0.000 352.270 4.000 ;
    END
  END wbs_adr_i[13]
  PIN wbs_adr_i[14]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 373.610 0.000 373.890 4.000 ;
    END
  END wbs_adr_i[14]
  PIN wbs_adr_i[15]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 394.770 0.000 395.050 4.000 ;
    END
  END wbs_adr_i[15]
  PIN wbs_adr_i[16]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 416.390 0.000 416.670 4.000 ;
    END
  END wbs_adr_i[16]
  PIN wbs_adr_i[17]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 437.550 0.000 437.830 4.000 ;
    END
  END wbs_adr_i[17]
  PIN wbs_adr_i[18]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 459.170 0.000 459.450 4.000 ;
    END
  END wbs_adr_i[18]
  PIN wbs_adr_i[19]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 480.330 0.000 480.610 4.000 ;
    END
  END wbs_adr_i[19]
  PIN wbs_adr_i[1]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 74.150 0.000 74.430 4.000 ;
    END
  END wbs_adr_i[1]
  PIN wbs_adr_i[20]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 501.950 0.000 502.230 4.000 ;
    END
  END wbs_adr_i[20]
  PIN wbs_adr_i[21]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 523.110 0.000 523.390 4.000 ;
    END
  END wbs_adr_i[21]
  PIN wbs_adr_i[22]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 544.270 0.000 544.550 4.000 ;
    END
  END wbs_adr_i[22]
  PIN wbs_adr_i[23]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 565.890 0.000 566.170 4.000 ;
    END
  END wbs_adr_i[23]
  PIN wbs_adr_i[24]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 587.050 0.000 587.330 4.000 ;
    END
  END wbs_adr_i[24]
  PIN wbs_adr_i[25]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 608.670 0.000 608.950 4.000 ;
    END
  END wbs_adr_i[25]
  PIN wbs_adr_i[26]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 629.830 0.000 630.110 4.000 ;
    END
  END wbs_adr_i[26]
  PIN wbs_adr_i[27]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 651.450 0.000 651.730 4.000 ;
    END
  END wbs_adr_i[27]
  PIN wbs_adr_i[28]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 672.610 0.000 672.890 4.000 ;
    END
  END wbs_adr_i[28]
  PIN wbs_adr_i[29]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 694.230 0.000 694.510 4.000 ;
    END
  END wbs_adr_i[29]
  PIN wbs_adr_i[2]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 102.670 0.000 102.950 4.000 ;
    END
  END wbs_adr_i[2]
  PIN wbs_adr_i[30]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 715.390 0.000 715.670 4.000 ;
    END
  END wbs_adr_i[30]
  PIN wbs_adr_i[31]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 737.010 0.000 737.290 4.000 ;
    END
  END wbs_adr_i[31]
  PIN wbs_adr_i[3]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 131.190 0.000 131.470 4.000 ;
    END
  END wbs_adr_i[3]
  PIN wbs_adr_i[4]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 159.710 0.000 159.990 4.000 ;
    END
  END wbs_adr_i[4]
  PIN wbs_adr_i[5]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 181.330 0.000 181.610 4.000 ;
    END
  END wbs_adr_i[5]
  PIN wbs_adr_i[6]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 202.490 0.000 202.770 4.000 ;
    END
  END wbs_adr_i[6]
  PIN wbs_adr_i[7]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 224.110 0.000 224.390 4.000 ;
    END
  END wbs_adr_i[7]
  PIN wbs_adr_i[8]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 245.270 0.000 245.550 4.000 ;
    END
  END wbs_adr_i[8]
  PIN wbs_adr_i[9]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 266.430 0.000 266.710 4.000 ;
    END
  END wbs_adr_i[9]
  PIN wbs_cyc_i
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 24.470 0.000 24.750 4.000 ;
    END
  END wbs_cyc_i
  PIN wbs_dat_i[0]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 52.990 0.000 53.270 4.000 ;
    END
  END wbs_dat_i[0]
  PIN wbs_dat_i[10]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 294.950 0.000 295.230 4.000 ;
    END
  END wbs_dat_i[10]
  PIN wbs_dat_i[11]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 316.570 0.000 316.850 4.000 ;
    END
  END wbs_dat_i[11]
  PIN wbs_dat_i[12]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 337.730 0.000 338.010 4.000 ;
    END
  END wbs_dat_i[12]
  PIN wbs_dat_i[13]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 359.350 0.000 359.630 4.000 ;
    END
  END wbs_dat_i[13]
  PIN wbs_dat_i[14]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 380.510 0.000 380.790 4.000 ;
    END
  END wbs_dat_i[14]
  PIN wbs_dat_i[15]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 402.130 0.000 402.410 4.000 ;
    END
  END wbs_dat_i[15]
  PIN wbs_dat_i[16]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 423.290 0.000 423.570 4.000 ;
    END
  END wbs_dat_i[16]
  PIN wbs_dat_i[17]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 444.910 0.000 445.190 4.000 ;
    END
  END wbs_dat_i[17]
  PIN wbs_dat_i[18]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 466.070 0.000 466.350 4.000 ;
    END
  END wbs_dat_i[18]
  PIN wbs_dat_i[19]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 487.690 0.000 487.970 4.000 ;
    END
  END wbs_dat_i[19]
  PIN wbs_dat_i[1]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 81.510 0.000 81.790 4.000 ;
    END
  END wbs_dat_i[1]
  PIN wbs_dat_i[20]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 508.850 0.000 509.130 4.000 ;
    END
  END wbs_dat_i[20]
  PIN wbs_dat_i[21]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 530.010 0.000 530.290 4.000 ;
    END
  END wbs_dat_i[21]
  PIN wbs_dat_i[22]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 551.630 0.000 551.910 4.000 ;
    END
  END wbs_dat_i[22]
  PIN wbs_dat_i[23]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 572.790 0.000 573.070 4.000 ;
    END
  END wbs_dat_i[23]
  PIN wbs_dat_i[24]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 594.410 0.000 594.690 4.000 ;
    END
  END wbs_dat_i[24]
  PIN wbs_dat_i[25]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 615.570 0.000 615.850 4.000 ;
    END
  END wbs_dat_i[25]
  PIN wbs_dat_i[26]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 637.190 0.000 637.470 4.000 ;
    END
  END wbs_dat_i[26]
  PIN wbs_dat_i[27]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 658.350 0.000 658.630 4.000 ;
    END
  END wbs_dat_i[27]
  PIN wbs_dat_i[28]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 679.970 0.000 680.250 4.000 ;
    END
  END wbs_dat_i[28]
  PIN wbs_dat_i[29]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 701.130 0.000 701.410 4.000 ;
    END
  END wbs_dat_i[29]
  PIN wbs_dat_i[2]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 110.030 0.000 110.310 4.000 ;
    END
  END wbs_dat_i[2]
  PIN wbs_dat_i[30]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 722.750 0.000 723.030 4.000 ;
    END
  END wbs_dat_i[30]
  PIN wbs_dat_i[31]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 743.910 0.000 744.190 4.000 ;
    END
  END wbs_dat_i[31]
  PIN wbs_dat_i[3]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 138.550 0.000 138.830 4.000 ;
    END
  END wbs_dat_i[3]
  PIN wbs_dat_i[4]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 167.070 0.000 167.350 4.000 ;
    END
  END wbs_dat_i[4]
  PIN wbs_dat_i[5]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 188.230 0.000 188.510 4.000 ;
    END
  END wbs_dat_i[5]
  PIN wbs_dat_i[6]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 209.850 0.000 210.130 4.000 ;
    END
  END wbs_dat_i[6]
  PIN wbs_dat_i[7]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 231.010 0.000 231.290 4.000 ;
    END
  END wbs_dat_i[7]
  PIN wbs_dat_i[8]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 252.630 0.000 252.910 4.000 ;
    END
  END wbs_dat_i[8]
  PIN wbs_dat_i[9]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 273.790 0.000 274.070 4.000 ;
    END
  END wbs_dat_i[9]
  PIN wbs_dat_o[0]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 59.890 0.000 60.170 4.000 ;
    END
  END wbs_dat_o[0]
  PIN wbs_dat_o[10]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 302.310 0.000 302.590 4.000 ;
    END
  END wbs_dat_o[10]
  PIN wbs_dat_o[11]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 323.470 0.000 323.750 4.000 ;
    END
  END wbs_dat_o[11]
  PIN wbs_dat_o[12]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 345.090 0.000 345.370 4.000 ;
    END
  END wbs_dat_o[12]
  PIN wbs_dat_o[13]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 366.250 0.000 366.530 4.000 ;
    END
  END wbs_dat_o[13]
  PIN wbs_dat_o[14]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 387.870 0.000 388.150 4.000 ;
    END
  END wbs_dat_o[14]
  PIN wbs_dat_o[15]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 409.030 0.000 409.310 4.000 ;
    END
  END wbs_dat_o[15]
  PIN wbs_dat_o[16]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 430.650 0.000 430.930 4.000 ;
    END
  END wbs_dat_o[16]
  PIN wbs_dat_o[17]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 451.810 0.000 452.090 4.000 ;
    END
  END wbs_dat_o[17]
  PIN wbs_dat_o[18]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 473.430 0.000 473.710 4.000 ;
    END
  END wbs_dat_o[18]
  PIN wbs_dat_o[19]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 494.590 0.000 494.870 4.000 ;
    END
  END wbs_dat_o[19]
  PIN wbs_dat_o[1]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 88.410 0.000 88.690 4.000 ;
    END
  END wbs_dat_o[1]
  PIN wbs_dat_o[20]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 515.750 0.000 516.030 4.000 ;
    END
  END wbs_dat_o[20]
  PIN wbs_dat_o[21]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 537.370 0.000 537.650 4.000 ;
    END
  END wbs_dat_o[21]
  PIN wbs_dat_o[22]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 558.530 0.000 558.810 4.000 ;
    END
  END wbs_dat_o[22]
  PIN wbs_dat_o[23]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 580.150 0.000 580.430 4.000 ;
    END
  END wbs_dat_o[23]
  PIN wbs_dat_o[24]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 601.310 0.000 601.590 4.000 ;
    END
  END wbs_dat_o[24]
  PIN wbs_dat_o[25]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 622.930 0.000 623.210 4.000 ;
    END
  END wbs_dat_o[25]
  PIN wbs_dat_o[26]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 644.090 0.000 644.370 4.000 ;
    END
  END wbs_dat_o[26]
  PIN wbs_dat_o[27]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 665.710 0.000 665.990 4.000 ;
    END
  END wbs_dat_o[27]
  PIN wbs_dat_o[28]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 686.870 0.000 687.150 4.000 ;
    END
  END wbs_dat_o[28]
  PIN wbs_dat_o[29]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 708.490 0.000 708.770 4.000 ;
    END
  END wbs_dat_o[29]
  PIN wbs_dat_o[2]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 116.930 0.000 117.210 4.000 ;
    END
  END wbs_dat_o[2]
  PIN wbs_dat_o[30]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 729.650 0.000 729.930 4.000 ;
    END
  END wbs_dat_o[30]
  PIN wbs_dat_o[31]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 751.270 0.000 751.550 4.000 ;
    END
  END wbs_dat_o[31]
  PIN wbs_dat_o[3]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 145.450 0.000 145.730 4.000 ;
    END
  END wbs_dat_o[3]
  PIN wbs_dat_o[4]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 173.970 0.000 174.250 4.000 ;
    END
  END wbs_dat_o[4]
  PIN wbs_dat_o[5]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 195.590 0.000 195.870 4.000 ;
    END
  END wbs_dat_o[5]
  PIN wbs_dat_o[6]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 216.750 0.000 217.030 4.000 ;
    END
  END wbs_dat_o[6]
  PIN wbs_dat_o[7]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 238.370 0.000 238.650 4.000 ;
    END
  END wbs_dat_o[7]
  PIN wbs_dat_o[8]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 259.530 0.000 259.810 4.000 ;
    END
  END wbs_dat_o[8]
  PIN wbs_dat_o[9]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 280.690 0.000 280.970 4.000 ;
    END
  END wbs_dat_o[9]
  PIN wbs_sel_i[0]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 67.250 0.000 67.530 4.000 ;
    END
  END wbs_sel_i[0]
  PIN wbs_sel_i[1]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 95.770 0.000 96.050 4.000 ;
    END
  END wbs_sel_i[1]
  PIN wbs_sel_i[2]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 124.290 0.000 124.570 4.000 ;
    END
  END wbs_sel_i[2]
  PIN wbs_sel_i[3]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 152.810 0.000 153.090 4.000 ;
    END
  END wbs_sel_i[3]
  PIN wbs_stb_i
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 31.370 0.000 31.650 4.000 ;
    END
  END wbs_stb_i
  PIN wbs_we_i
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 38.730 0.000 39.010 4.000 ;
    END
  END wbs_we_i
  OBS
      LAYER li1 ;
        RECT 5.520 10.795 995.755 995.605 ;
      LAYER met1 ;
        RECT 5.520 2.420 996.750 997.180 ;
      LAYER met2 ;
        RECT 3.410 1003.560 8.550 1003.840 ;
        RECT 9.390 1003.560 14.990 1003.840 ;
        RECT 15.830 1003.560 20.970 1003.840 ;
        RECT 21.810 1003.560 27.410 1003.840 ;
        RECT 28.250 1003.560 33.850 1003.840 ;
        RECT 34.690 1003.560 39.830 1003.840 ;
        RECT 40.670 1003.560 46.270 1003.840 ;
        RECT 47.110 1003.560 52.710 1003.840 ;
        RECT 53.550 1003.560 58.690 1003.840 ;
        RECT 59.530 1003.560 65.130 1003.840 ;
        RECT 65.970 1003.560 71.110 1003.840 ;
        RECT 71.950 1003.560 77.550 1003.840 ;
        RECT 78.390 1003.560 83.990 1003.840 ;
        RECT 84.830 1003.560 89.970 1003.840 ;
        RECT 90.810 1003.560 96.410 1003.840 ;
        RECT 97.250 1003.560 102.850 1003.840 ;
        RECT 103.690 1003.560 108.830 1003.840 ;
        RECT 109.670 1003.560 115.270 1003.840 ;
        RECT 116.110 1003.560 121.710 1003.840 ;
        RECT 122.550 1003.560 127.690 1003.840 ;
        RECT 128.530 1003.560 134.130 1003.840 ;
        RECT 134.970 1003.560 140.110 1003.840 ;
        RECT 140.950 1003.560 146.550 1003.840 ;
        RECT 147.390 1003.560 152.990 1003.840 ;
        RECT 153.830 1003.560 158.970 1003.840 ;
        RECT 159.810 1003.560 165.410 1003.840 ;
        RECT 166.250 1003.560 171.850 1003.840 ;
        RECT 172.690 1003.560 177.830 1003.840 ;
        RECT 178.670 1003.560 184.270 1003.840 ;
        RECT 185.110 1003.560 190.710 1003.840 ;
        RECT 191.550 1003.560 196.690 1003.840 ;
        RECT 197.530 1003.560 203.130 1003.840 ;
        RECT 203.970 1003.560 209.110 1003.840 ;
        RECT 209.950 1003.560 215.550 1003.840 ;
        RECT 216.390 1003.560 221.990 1003.840 ;
        RECT 222.830 1003.560 227.970 1003.840 ;
        RECT 228.810 1003.560 234.410 1003.840 ;
        RECT 235.250 1003.560 240.850 1003.840 ;
        RECT 241.690 1003.560 246.830 1003.840 ;
        RECT 247.670 1003.560 253.270 1003.840 ;
        RECT 254.110 1003.560 259.710 1003.840 ;
        RECT 260.550 1003.560 265.690 1003.840 ;
        RECT 266.530 1003.560 272.130 1003.840 ;
        RECT 272.970 1003.560 278.110 1003.840 ;
        RECT 278.950 1003.560 284.550 1003.840 ;
        RECT 285.390 1003.560 290.990 1003.840 ;
        RECT 291.830 1003.560 296.970 1003.840 ;
        RECT 297.810 1003.560 303.410 1003.840 ;
        RECT 304.250 1003.560 309.850 1003.840 ;
        RECT 310.690 1003.560 315.830 1003.840 ;
        RECT 316.670 1003.560 322.270 1003.840 ;
        RECT 323.110 1003.560 328.710 1003.840 ;
        RECT 329.550 1003.560 334.690 1003.840 ;
        RECT 335.530 1003.560 341.130 1003.840 ;
        RECT 341.970 1003.560 347.110 1003.840 ;
        RECT 347.950 1003.560 353.550 1003.840 ;
        RECT 354.390 1003.560 359.990 1003.840 ;
        RECT 360.830 1003.560 365.970 1003.840 ;
        RECT 366.810 1003.560 372.410 1003.840 ;
        RECT 373.250 1003.560 378.850 1003.840 ;
        RECT 379.690 1003.560 384.830 1003.840 ;
        RECT 385.670 1003.560 391.270 1003.840 ;
        RECT 392.110 1003.560 397.710 1003.840 ;
        RECT 398.550 1003.560 403.690 1003.840 ;
        RECT 404.530 1003.560 410.130 1003.840 ;
        RECT 410.970 1003.560 416.110 1003.840 ;
        RECT 416.950 1003.560 422.550 1003.840 ;
        RECT 423.390 1003.560 428.990 1003.840 ;
        RECT 429.830 1003.560 434.970 1003.840 ;
        RECT 435.810 1003.560 441.410 1003.840 ;
        RECT 442.250 1003.560 447.850 1003.840 ;
        RECT 448.690 1003.560 453.830 1003.840 ;
        RECT 454.670 1003.560 460.270 1003.840 ;
        RECT 461.110 1003.560 466.710 1003.840 ;
        RECT 467.550 1003.560 472.690 1003.840 ;
        RECT 473.530 1003.560 479.130 1003.840 ;
        RECT 479.970 1003.560 485.110 1003.840 ;
        RECT 485.950 1003.560 491.550 1003.840 ;
        RECT 492.390 1003.560 497.990 1003.840 ;
        RECT 498.830 1003.560 503.970 1003.840 ;
        RECT 504.810 1003.560 510.410 1003.840 ;
        RECT 511.250 1003.560 516.850 1003.840 ;
        RECT 517.690 1003.560 522.830 1003.840 ;
        RECT 523.670 1003.560 529.270 1003.840 ;
        RECT 530.110 1003.560 535.250 1003.840 ;
        RECT 536.090 1003.560 541.690 1003.840 ;
        RECT 542.530 1003.560 548.130 1003.840 ;
        RECT 548.970 1003.560 554.110 1003.840 ;
        RECT 554.950 1003.560 560.550 1003.840 ;
        RECT 561.390 1003.560 566.990 1003.840 ;
        RECT 567.830 1003.560 572.970 1003.840 ;
        RECT 573.810 1003.560 579.410 1003.840 ;
        RECT 580.250 1003.560 585.850 1003.840 ;
        RECT 586.690 1003.560 591.830 1003.840 ;
        RECT 592.670 1003.560 598.270 1003.840 ;
        RECT 599.110 1003.560 604.250 1003.840 ;
        RECT 605.090 1003.560 610.690 1003.840 ;
        RECT 611.530 1003.560 617.130 1003.840 ;
        RECT 617.970 1003.560 623.110 1003.840 ;
        RECT 623.950 1003.560 629.550 1003.840 ;
        RECT 630.390 1003.560 635.990 1003.840 ;
        RECT 636.830 1003.560 641.970 1003.840 ;
        RECT 642.810 1003.560 648.410 1003.840 ;
        RECT 649.250 1003.560 654.850 1003.840 ;
        RECT 655.690 1003.560 660.830 1003.840 ;
        RECT 661.670 1003.560 667.270 1003.840 ;
        RECT 668.110 1003.560 673.250 1003.840 ;
        RECT 674.090 1003.560 679.690 1003.840 ;
        RECT 680.530 1003.560 686.130 1003.840 ;
        RECT 686.970 1003.560 692.110 1003.840 ;
        RECT 692.950 1003.560 698.550 1003.840 ;
        RECT 699.390 1003.560 704.990 1003.840 ;
        RECT 705.830 1003.560 710.970 1003.840 ;
        RECT 711.810 1003.560 717.410 1003.840 ;
        RECT 718.250 1003.560 723.850 1003.840 ;
        RECT 724.690 1003.560 729.830 1003.840 ;
        RECT 730.670 1003.560 736.270 1003.840 ;
        RECT 737.110 1003.560 742.250 1003.840 ;
        RECT 743.090 1003.560 748.690 1003.840 ;
        RECT 749.530 1003.560 755.130 1003.840 ;
        RECT 755.970 1003.560 761.110 1003.840 ;
        RECT 761.950 1003.560 767.550 1003.840 ;
        RECT 768.390 1003.560 773.990 1003.840 ;
        RECT 774.830 1003.560 779.970 1003.840 ;
        RECT 780.810 1003.560 786.410 1003.840 ;
        RECT 787.250 1003.560 792.850 1003.840 ;
        RECT 793.690 1003.560 798.830 1003.840 ;
        RECT 799.670 1003.560 805.270 1003.840 ;
        RECT 806.110 1003.560 811.250 1003.840 ;
        RECT 812.090 1003.560 817.690 1003.840 ;
        RECT 818.530 1003.560 824.130 1003.840 ;
        RECT 824.970 1003.560 830.110 1003.840 ;
        RECT 830.950 1003.560 836.550 1003.840 ;
        RECT 837.390 1003.560 842.990 1003.840 ;
        RECT 843.830 1003.560 848.970 1003.840 ;
        RECT 849.810 1003.560 855.410 1003.840 ;
        RECT 856.250 1003.560 861.850 1003.840 ;
        RECT 862.690 1003.560 867.830 1003.840 ;
        RECT 868.670 1003.560 874.270 1003.840 ;
        RECT 875.110 1003.560 880.250 1003.840 ;
        RECT 881.090 1003.560 886.690 1003.840 ;
        RECT 887.530 1003.560 893.130 1003.840 ;
        RECT 893.970 1003.560 899.110 1003.840 ;
        RECT 899.950 1003.560 905.550 1003.840 ;
        RECT 906.390 1003.560 911.990 1003.840 ;
        RECT 912.830 1003.560 917.970 1003.840 ;
        RECT 918.810 1003.560 924.410 1003.840 ;
        RECT 925.250 1003.560 930.850 1003.840 ;
        RECT 931.690 1003.560 936.830 1003.840 ;
        RECT 937.670 1003.560 943.270 1003.840 ;
        RECT 944.110 1003.560 949.250 1003.840 ;
        RECT 950.090 1003.560 955.690 1003.840 ;
        RECT 956.530 1003.560 962.130 1003.840 ;
        RECT 962.970 1003.560 968.110 1003.840 ;
        RECT 968.950 1003.560 974.550 1003.840 ;
        RECT 975.390 1003.560 980.990 1003.840 ;
        RECT 981.830 1003.560 986.970 1003.840 ;
        RECT 987.810 1003.560 993.410 1003.840 ;
        RECT 994.250 1003.560 996.720 1003.840 ;
        RECT 3.380 4.280 996.720 1003.560 ;
        RECT 3.870 0.155 9.930 4.280 ;
        RECT 10.770 0.155 16.830 4.280 ;
        RECT 17.670 0.155 24.190 4.280 ;
        RECT 25.030 0.155 31.090 4.280 ;
        RECT 31.930 0.155 38.450 4.280 ;
        RECT 39.290 0.155 45.350 4.280 ;
        RECT 46.190 0.155 52.710 4.280 ;
        RECT 53.550 0.155 59.610 4.280 ;
        RECT 60.450 0.155 66.970 4.280 ;
        RECT 67.810 0.155 73.870 4.280 ;
        RECT 74.710 0.155 81.230 4.280 ;
        RECT 82.070 0.155 88.130 4.280 ;
        RECT 88.970 0.155 95.490 4.280 ;
        RECT 96.330 0.155 102.390 4.280 ;
        RECT 103.230 0.155 109.750 4.280 ;
        RECT 110.590 0.155 116.650 4.280 ;
        RECT 117.490 0.155 124.010 4.280 ;
        RECT 124.850 0.155 130.910 4.280 ;
        RECT 131.750 0.155 138.270 4.280 ;
        RECT 139.110 0.155 145.170 4.280 ;
        RECT 146.010 0.155 152.530 4.280 ;
        RECT 153.370 0.155 159.430 4.280 ;
        RECT 160.270 0.155 166.790 4.280 ;
        RECT 167.630 0.155 173.690 4.280 ;
        RECT 174.530 0.155 181.050 4.280 ;
        RECT 181.890 0.155 187.950 4.280 ;
        RECT 188.790 0.155 195.310 4.280 ;
        RECT 196.150 0.155 202.210 4.280 ;
        RECT 203.050 0.155 209.570 4.280 ;
        RECT 210.410 0.155 216.470 4.280 ;
        RECT 217.310 0.155 223.830 4.280 ;
        RECT 224.670 0.155 230.730 4.280 ;
        RECT 231.570 0.155 238.090 4.280 ;
        RECT 238.930 0.155 244.990 4.280 ;
        RECT 245.830 0.155 252.350 4.280 ;
        RECT 253.190 0.155 259.250 4.280 ;
        RECT 260.090 0.155 266.150 4.280 ;
        RECT 266.990 0.155 273.510 4.280 ;
        RECT 274.350 0.155 280.410 4.280 ;
        RECT 281.250 0.155 287.770 4.280 ;
        RECT 288.610 0.155 294.670 4.280 ;
        RECT 295.510 0.155 302.030 4.280 ;
        RECT 302.870 0.155 308.930 4.280 ;
        RECT 309.770 0.155 316.290 4.280 ;
        RECT 317.130 0.155 323.190 4.280 ;
        RECT 324.030 0.155 330.550 4.280 ;
        RECT 331.390 0.155 337.450 4.280 ;
        RECT 338.290 0.155 344.810 4.280 ;
        RECT 345.650 0.155 351.710 4.280 ;
        RECT 352.550 0.155 359.070 4.280 ;
        RECT 359.910 0.155 365.970 4.280 ;
        RECT 366.810 0.155 373.330 4.280 ;
        RECT 374.170 0.155 380.230 4.280 ;
        RECT 381.070 0.155 387.590 4.280 ;
        RECT 388.430 0.155 394.490 4.280 ;
        RECT 395.330 0.155 401.850 4.280 ;
        RECT 402.690 0.155 408.750 4.280 ;
        RECT 409.590 0.155 416.110 4.280 ;
        RECT 416.950 0.155 423.010 4.280 ;
        RECT 423.850 0.155 430.370 4.280 ;
        RECT 431.210 0.155 437.270 4.280 ;
        RECT 438.110 0.155 444.630 4.280 ;
        RECT 445.470 0.155 451.530 4.280 ;
        RECT 452.370 0.155 458.890 4.280 ;
        RECT 459.730 0.155 465.790 4.280 ;
        RECT 466.630 0.155 473.150 4.280 ;
        RECT 473.990 0.155 480.050 4.280 ;
        RECT 480.890 0.155 487.410 4.280 ;
        RECT 488.250 0.155 494.310 4.280 ;
        RECT 495.150 0.155 501.670 4.280 ;
        RECT 502.510 0.155 508.570 4.280 ;
        RECT 509.410 0.155 515.470 4.280 ;
        RECT 516.310 0.155 522.830 4.280 ;
        RECT 523.670 0.155 529.730 4.280 ;
        RECT 530.570 0.155 537.090 4.280 ;
        RECT 537.930 0.155 543.990 4.280 ;
        RECT 544.830 0.155 551.350 4.280 ;
        RECT 552.190 0.155 558.250 4.280 ;
        RECT 559.090 0.155 565.610 4.280 ;
        RECT 566.450 0.155 572.510 4.280 ;
        RECT 573.350 0.155 579.870 4.280 ;
        RECT 580.710 0.155 586.770 4.280 ;
        RECT 587.610 0.155 594.130 4.280 ;
        RECT 594.970 0.155 601.030 4.280 ;
        RECT 601.870 0.155 608.390 4.280 ;
        RECT 609.230 0.155 615.290 4.280 ;
        RECT 616.130 0.155 622.650 4.280 ;
        RECT 623.490 0.155 629.550 4.280 ;
        RECT 630.390 0.155 636.910 4.280 ;
        RECT 637.750 0.155 643.810 4.280 ;
        RECT 644.650 0.155 651.170 4.280 ;
        RECT 652.010 0.155 658.070 4.280 ;
        RECT 658.910 0.155 665.430 4.280 ;
        RECT 666.270 0.155 672.330 4.280 ;
        RECT 673.170 0.155 679.690 4.280 ;
        RECT 680.530 0.155 686.590 4.280 ;
        RECT 687.430 0.155 693.950 4.280 ;
        RECT 694.790 0.155 700.850 4.280 ;
        RECT 701.690 0.155 708.210 4.280 ;
        RECT 709.050 0.155 715.110 4.280 ;
        RECT 715.950 0.155 722.470 4.280 ;
        RECT 723.310 0.155 729.370 4.280 ;
        RECT 730.210 0.155 736.730 4.280 ;
        RECT 737.570 0.155 743.630 4.280 ;
        RECT 744.470 0.155 750.990 4.280 ;
        RECT 751.830 0.155 757.890 4.280 ;
        RECT 758.730 0.155 764.790 4.280 ;
        RECT 765.630 0.155 772.150 4.280 ;
        RECT 772.990 0.155 779.050 4.280 ;
        RECT 779.890 0.155 786.410 4.280 ;
        RECT 787.250 0.155 793.310 4.280 ;
        RECT 794.150 0.155 800.670 4.280 ;
        RECT 801.510 0.155 807.570 4.280 ;
        RECT 808.410 0.155 814.930 4.280 ;
        RECT 815.770 0.155 821.830 4.280 ;
        RECT 822.670 0.155 829.190 4.280 ;
        RECT 830.030 0.155 836.090 4.280 ;
        RECT 836.930 0.155 843.450 4.280 ;
        RECT 844.290 0.155 850.350 4.280 ;
        RECT 851.190 0.155 857.710 4.280 ;
        RECT 858.550 0.155 864.610 4.280 ;
        RECT 865.450 0.155 871.970 4.280 ;
        RECT 872.810 0.155 878.870 4.280 ;
        RECT 879.710 0.155 886.230 4.280 ;
        RECT 887.070 0.155 893.130 4.280 ;
        RECT 893.970 0.155 900.490 4.280 ;
        RECT 901.330 0.155 907.390 4.280 ;
        RECT 908.230 0.155 914.750 4.280 ;
        RECT 915.590 0.155 921.650 4.280 ;
        RECT 922.490 0.155 929.010 4.280 ;
        RECT 929.850 0.155 935.910 4.280 ;
        RECT 936.750 0.155 943.270 4.280 ;
        RECT 944.110 0.155 950.170 4.280 ;
        RECT 951.010 0.155 957.530 4.280 ;
        RECT 958.370 0.155 964.430 4.280 ;
        RECT 965.270 0.155 971.790 4.280 ;
        RECT 972.630 0.155 978.690 4.280 ;
        RECT 979.530 0.155 986.050 4.280 ;
        RECT 986.890 0.155 992.950 4.280 ;
        RECT 993.790 0.155 996.720 4.280 ;
      LAYER met3 ;
        RECT 3.745 997.240 996.295 998.065 ;
        RECT 4.400 995.840 996.295 997.240 ;
        RECT 3.745 995.200 996.295 995.840 ;
        RECT 3.745 993.800 992.720 995.200 ;
        RECT 3.745 975.480 996.295 993.800 ;
        RECT 4.400 974.080 996.295 975.480 ;
        RECT 3.745 968.680 996.295 974.080 ;
        RECT 3.745 967.280 992.720 968.680 ;
        RECT 3.745 953.720 996.295 967.280 ;
        RECT 4.400 952.320 996.295 953.720 ;
        RECT 3.745 942.160 996.295 952.320 ;
        RECT 3.745 940.760 992.720 942.160 ;
        RECT 3.745 931.960 996.295 940.760 ;
        RECT 4.400 930.560 996.295 931.960 ;
        RECT 3.745 915.640 996.295 930.560 ;
        RECT 3.745 914.240 992.720 915.640 ;
        RECT 3.745 909.520 996.295 914.240 ;
        RECT 4.400 908.120 996.295 909.520 ;
        RECT 3.745 889.120 996.295 908.120 ;
        RECT 3.745 887.760 992.720 889.120 ;
        RECT 4.400 887.720 992.720 887.760 ;
        RECT 4.400 886.360 996.295 887.720 ;
        RECT 3.745 866.000 996.295 886.360 ;
        RECT 4.400 864.600 996.295 866.000 ;
        RECT 3.745 862.600 996.295 864.600 ;
        RECT 3.745 861.200 992.720 862.600 ;
        RECT 3.745 844.240 996.295 861.200 ;
        RECT 4.400 842.840 996.295 844.240 ;
        RECT 3.745 836.080 996.295 842.840 ;
        RECT 3.745 834.680 992.720 836.080 ;
        RECT 3.745 822.480 996.295 834.680 ;
        RECT 4.400 821.080 996.295 822.480 ;
        RECT 3.745 809.560 996.295 821.080 ;
        RECT 3.745 808.160 992.720 809.560 ;
        RECT 3.745 800.040 996.295 808.160 ;
        RECT 4.400 798.640 996.295 800.040 ;
        RECT 3.745 783.040 996.295 798.640 ;
        RECT 3.745 781.640 992.720 783.040 ;
        RECT 3.745 778.280 996.295 781.640 ;
        RECT 4.400 776.880 996.295 778.280 ;
        RECT 3.745 756.520 996.295 776.880 ;
        RECT 4.400 755.120 992.720 756.520 ;
        RECT 3.745 734.760 996.295 755.120 ;
        RECT 4.400 733.360 996.295 734.760 ;
        RECT 3.745 730.000 996.295 733.360 ;
        RECT 3.745 728.600 992.720 730.000 ;
        RECT 3.745 712.320 996.295 728.600 ;
        RECT 4.400 710.920 996.295 712.320 ;
        RECT 3.745 703.480 996.295 710.920 ;
        RECT 3.745 702.080 992.720 703.480 ;
        RECT 3.745 690.560 996.295 702.080 ;
        RECT 4.400 689.160 996.295 690.560 ;
        RECT 3.745 676.960 996.295 689.160 ;
        RECT 3.745 675.560 992.720 676.960 ;
        RECT 3.745 668.800 996.295 675.560 ;
        RECT 4.400 667.400 996.295 668.800 ;
        RECT 3.745 650.440 996.295 667.400 ;
        RECT 3.745 649.040 992.720 650.440 ;
        RECT 3.745 647.040 996.295 649.040 ;
        RECT 4.400 645.640 996.295 647.040 ;
        RECT 3.745 625.280 996.295 645.640 ;
        RECT 4.400 623.920 996.295 625.280 ;
        RECT 4.400 623.880 992.720 623.920 ;
        RECT 3.745 622.520 992.720 623.880 ;
        RECT 3.745 602.840 996.295 622.520 ;
        RECT 4.400 601.440 996.295 602.840 ;
        RECT 3.745 597.400 996.295 601.440 ;
        RECT 3.745 596.000 992.720 597.400 ;
        RECT 3.745 581.080 996.295 596.000 ;
        RECT 4.400 579.680 996.295 581.080 ;
        RECT 3.745 570.880 996.295 579.680 ;
        RECT 3.745 569.480 992.720 570.880 ;
        RECT 3.745 559.320 996.295 569.480 ;
        RECT 4.400 557.920 996.295 559.320 ;
        RECT 3.745 544.360 996.295 557.920 ;
        RECT 3.745 542.960 992.720 544.360 ;
        RECT 3.745 537.560 996.295 542.960 ;
        RECT 4.400 536.160 996.295 537.560 ;
        RECT 3.745 517.840 996.295 536.160 ;
        RECT 3.745 516.440 992.720 517.840 ;
        RECT 3.745 515.800 996.295 516.440 ;
        RECT 4.400 514.400 996.295 515.800 ;
        RECT 3.745 493.360 996.295 514.400 ;
        RECT 4.400 491.960 996.295 493.360 ;
        RECT 3.745 491.320 996.295 491.960 ;
        RECT 3.745 489.920 992.720 491.320 ;
        RECT 3.745 471.600 996.295 489.920 ;
        RECT 4.400 470.200 996.295 471.600 ;
        RECT 3.745 464.800 996.295 470.200 ;
        RECT 3.745 463.400 992.720 464.800 ;
        RECT 3.745 449.840 996.295 463.400 ;
        RECT 4.400 448.440 996.295 449.840 ;
        RECT 3.745 438.280 996.295 448.440 ;
        RECT 3.745 436.880 992.720 438.280 ;
        RECT 3.745 428.080 996.295 436.880 ;
        RECT 4.400 426.680 996.295 428.080 ;
        RECT 3.745 411.760 996.295 426.680 ;
        RECT 3.745 410.360 992.720 411.760 ;
        RECT 3.745 405.640 996.295 410.360 ;
        RECT 4.400 404.240 996.295 405.640 ;
        RECT 3.745 385.240 996.295 404.240 ;
        RECT 3.745 383.880 992.720 385.240 ;
        RECT 4.400 383.840 992.720 383.880 ;
        RECT 4.400 382.480 996.295 383.840 ;
        RECT 3.745 362.120 996.295 382.480 ;
        RECT 4.400 360.720 996.295 362.120 ;
        RECT 3.745 358.720 996.295 360.720 ;
        RECT 3.745 357.320 992.720 358.720 ;
        RECT 3.745 340.360 996.295 357.320 ;
        RECT 4.400 338.960 996.295 340.360 ;
        RECT 3.745 332.200 996.295 338.960 ;
        RECT 3.745 330.800 992.720 332.200 ;
        RECT 3.745 318.600 996.295 330.800 ;
        RECT 4.400 317.200 996.295 318.600 ;
        RECT 3.745 305.680 996.295 317.200 ;
        RECT 3.745 304.280 992.720 305.680 ;
        RECT 3.745 296.160 996.295 304.280 ;
        RECT 4.400 294.760 996.295 296.160 ;
        RECT 3.745 279.160 996.295 294.760 ;
        RECT 3.745 277.760 992.720 279.160 ;
        RECT 3.745 274.400 996.295 277.760 ;
        RECT 4.400 273.000 996.295 274.400 ;
        RECT 3.745 252.640 996.295 273.000 ;
        RECT 4.400 251.240 992.720 252.640 ;
        RECT 3.745 230.880 996.295 251.240 ;
        RECT 4.400 229.480 996.295 230.880 ;
        RECT 3.745 226.120 996.295 229.480 ;
        RECT 3.745 224.720 992.720 226.120 ;
        RECT 3.745 208.440 996.295 224.720 ;
        RECT 4.400 207.040 996.295 208.440 ;
        RECT 3.745 199.600 996.295 207.040 ;
        RECT 3.745 198.200 992.720 199.600 ;
        RECT 3.745 186.680 996.295 198.200 ;
        RECT 4.400 185.280 996.295 186.680 ;
        RECT 3.745 173.080 996.295 185.280 ;
        RECT 3.745 171.680 992.720 173.080 ;
        RECT 3.745 164.920 996.295 171.680 ;
        RECT 4.400 163.520 996.295 164.920 ;
        RECT 3.745 146.560 996.295 163.520 ;
        RECT 3.745 145.160 992.720 146.560 ;
        RECT 3.745 143.160 996.295 145.160 ;
        RECT 4.400 141.760 996.295 143.160 ;
        RECT 3.745 121.400 996.295 141.760 ;
        RECT 4.400 120.040 996.295 121.400 ;
        RECT 4.400 120.000 992.720 120.040 ;
        RECT 3.745 118.640 992.720 120.000 ;
        RECT 3.745 98.960 996.295 118.640 ;
        RECT 4.400 97.560 996.295 98.960 ;
        RECT 3.745 93.520 996.295 97.560 ;
        RECT 3.745 92.120 992.720 93.520 ;
        RECT 3.745 77.200 996.295 92.120 ;
        RECT 4.400 75.800 996.295 77.200 ;
        RECT 3.745 67.000 996.295 75.800 ;
        RECT 3.745 65.600 992.720 67.000 ;
        RECT 3.745 55.440 996.295 65.600 ;
        RECT 4.400 54.040 996.295 55.440 ;
        RECT 3.745 40.480 996.295 54.040 ;
        RECT 3.745 39.080 992.720 40.480 ;
        RECT 3.745 33.680 996.295 39.080 ;
        RECT 4.400 32.280 996.295 33.680 ;
        RECT 3.745 13.960 996.295 32.280 ;
        RECT 3.745 12.560 992.720 13.960 ;
        RECT 3.745 11.920 996.295 12.560 ;
        RECT 4.400 10.520 996.295 11.920 ;
        RECT 3.745 0.175 996.295 10.520 ;
      LAYER met4 ;
        RECT 44.455 996.160 983.185 998.065 ;
        RECT 44.455 10.240 97.440 996.160 ;
        RECT 99.840 10.240 174.240 996.160 ;
        RECT 176.640 10.240 251.040 996.160 ;
        RECT 253.440 10.240 327.840 996.160 ;
        RECT 330.240 10.240 404.640 996.160 ;
        RECT 407.040 10.240 481.440 996.160 ;
        RECT 483.840 10.240 558.240 996.160 ;
        RECT 560.640 10.240 635.040 996.160 ;
        RECT 637.440 10.240 711.840 996.160 ;
        RECT 714.240 10.240 788.640 996.160 ;
        RECT 791.040 10.240 865.440 996.160 ;
        RECT 867.840 10.240 942.240 996.160 ;
        RECT 944.640 10.240 983.185 996.160 ;
        RECT 44.455 5.615 983.185 10.240 ;
  END
END user_proj
END LIBRARY

