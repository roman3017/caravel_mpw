VERSION 5.7 ;
  NOWIREEXTENSIONATPIN ON ;
  DIVIDERCHAR "/" ;
  BUSBITCHARS "[]" ;
MACRO user_proj
  CLASS BLOCK ;
  FOREIGN user_proj ;
  ORIGIN 0.000 0.000 ;
  SIZE 990.625 BY 1001.345 ;
  PIN clk_i
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 986.625 15.680 990.625 16.280 ;
    END
  END clk_i
  PIN i_dout0[0]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 731.490 997.345 731.770 1001.345 ;
    END
  END i_dout0[0]
  PIN i_dout0[10]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 818.890 0.000 819.170 4.000 ;
    END
  END i_dout0[10]
  PIN i_dout0[11]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 832.230 0.000 832.510 4.000 ;
    END
  END i_dout0[11]
  PIN i_dout0[12]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 845.110 0.000 845.390 4.000 ;
    END
  END i_dout0[12]
  PIN i_dout0[13]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 986.625 499.840 990.625 500.440 ;
    END
  END i_dout0[13]
  PIN i_dout0[14]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 579.400 4.000 580.000 ;
    END
  END i_dout0[14]
  PIN i_dout0[15]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 602.520 4.000 603.120 ;
    END
  END i_dout0[15]
  PIN i_dout0[16]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 884.670 997.345 884.950 1001.345 ;
    END
  END i_dout0[16]
  PIN i_dout0[17]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 877.310 0.000 877.590 4.000 ;
    END
  END i_dout0[17]
  PIN i_dout0[18]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 897.550 997.345 897.830 1001.345 ;
    END
  END i_dout0[18]
  PIN i_dout0[19]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 890.190 0.000 890.470 4.000 ;
    END
  END i_dout0[19]
  PIN i_dout0[1]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 986.625 144.880 990.625 145.480 ;
    END
  END i_dout0[1]
  PIN i_dout0[20]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 903.990 997.345 904.270 1001.345 ;
    END
  END i_dout0[20]
  PIN i_dout0[21]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 896.630 0.000 896.910 4.000 ;
    END
  END i_dout0[21]
  PIN i_dout0[22]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 852.760 4.000 853.360 ;
    END
  END i_dout0[22]
  PIN i_dout0[23]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 875.880 4.000 876.480 ;
    END
  END i_dout0[23]
  PIN i_dout0[24]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 898.320 4.000 898.920 ;
    END
  END i_dout0[24]
  PIN i_dout0[25]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 921.440 4.000 922.040 ;
    END
  END i_dout0[25]
  PIN i_dout0[26]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 967.930 997.345 968.210 1001.345 ;
    END
  END i_dout0[26]
  PIN i_dout0[27]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 922.850 0.000 923.130 4.000 ;
    END
  END i_dout0[27]
  PIN i_dout0[28]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 986.625 920.080 990.625 920.680 ;
    END
  END i_dout0[28]
  PIN i_dout0[29]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 980.810 997.345 981.090 1001.345 ;
    END
  END i_dout0[29]
  PIN i_dout0[2]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 215.600 4.000 216.200 ;
    END
  END i_dout0[2]
  PIN i_dout0[30]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 961.490 0.000 961.770 4.000 ;
    END
  END i_dout0[30]
  PIN i_dout0[31]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 986.625 984.680 990.625 985.280 ;
    END
  END i_dout0[31]
  PIN i_dout0[3]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 238.040 4.000 238.640 ;
    END
  END i_dout0[3]
  PIN i_dout0[4]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 306.720 4.000 307.320 ;
    END
  END i_dout0[4]
  PIN i_dout0[5]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 767.370 0.000 767.650 4.000 ;
    END
  END i_dout0[5]
  PIN i_dout0[6]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 986.625 338.680 990.625 339.280 ;
    END
  END i_dout0[6]
  PIN i_dout0[7]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 820.730 997.345 821.010 1001.345 ;
    END
  END i_dout0[7]
  PIN i_dout0[8]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 443.400 4.000 444.000 ;
    END
  END i_dout0[8]
  PIN i_dout0[9]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 511.400 4.000 512.000 ;
    END
  END i_dout0[9]
  PIN i_dout0_1[0]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 55.800 4.000 56.400 ;
    END
  END i_dout0_1[0]
  PIN i_dout0_1[10]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 852.930 997.345 853.210 1001.345 ;
    END
  END i_dout0_1[10]
  PIN i_dout0_1[11]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 825.330 0.000 825.610 4.000 ;
    END
  END i_dout0_1[11]
  PIN i_dout0_1[12]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 838.670 0.000 838.950 4.000 ;
    END
  END i_dout0_1[12]
  PIN i_dout0_1[13]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 533.840 4.000 534.440 ;
    END
  END i_dout0_1[13]
  PIN i_dout0_1[14]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 986.625 532.480 990.625 533.080 ;
    END
  END i_dout0_1[14]
  PIN i_dout0_1[15]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 878.230 997.345 878.510 1001.345 ;
    END
  END i_dout0_1[15]
  PIN i_dout0_1[16]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 624.960 4.000 625.560 ;
    END
  END i_dout0_1[16]
  PIN i_dout0_1[17]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 648.080 4.000 648.680 ;
    END
  END i_dout0_1[17]
  PIN i_dout0_1[18]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 986.625 661.680 990.625 662.280 ;
    END
  END i_dout0_1[18]
  PIN i_dout0_1[19]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 739.200 4.000 739.800 ;
    END
  END i_dout0_1[19]
  PIN i_dout0_1[1]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 146.920 4.000 147.520 ;
    END
  END i_dout0_1[1]
  PIN i_dout0_1[20]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 986.625 726.280 990.625 726.880 ;
    END
  END i_dout0_1[20]
  PIN i_dout0_1[21]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 807.200 4.000 807.800 ;
    END
  END i_dout0_1[21]
  PIN i_dout0_1[22]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 916.870 997.345 917.150 1001.345 ;
    END
  END i_dout0_1[22]
  PIN i_dout0_1[23]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 923.310 997.345 923.590 1001.345 ;
    END
  END i_dout0_1[23]
  PIN i_dout0_1[24]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 903.070 0.000 903.350 4.000 ;
    END
  END i_dout0_1[24]
  PIN i_dout0_1[25]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 948.610 997.345 948.890 1001.345 ;
    END
  END i_dout0_1[25]
  PIN i_dout0_1[26]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 943.880 4.000 944.480 ;
    END
  END i_dout0_1[26]
  PIN i_dout0_1[27]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 916.410 0.000 916.690 4.000 ;
    END
  END i_dout0_1[27]
  PIN i_dout0_1[28]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 935.730 0.000 936.010 4.000 ;
    END
  END i_dout0_1[28]
  PIN i_dout0_1[29]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 974.370 997.345 974.650 1001.345 ;
    END
  END i_dout0_1[29]
  PIN i_dout0_1[2]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 986.625 209.480 990.625 210.080 ;
    END
  END i_dout0_1[2]
  PIN i_dout0_1[30]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 955.050 0.000 955.330 4.000 ;
    END
  END i_dout0_1[30]
  PIN i_dout0_1[31]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 980.810 0.000 981.090 4.000 ;
    END
  END i_dout0_1[31]
  PIN i_dout0_1[3]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 748.050 0.000 748.330 4.000 ;
    END
  END i_dout0_1[3]
  PIN i_dout0_1[4]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 986.625 306.040 990.625 306.640 ;
    END
  END i_dout0_1[4]
  PIN i_dout0_1[5]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 795.430 997.345 795.710 1001.345 ;
    END
  END i_dout0_1[5]
  PIN i_dout0_1[6]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 397.840 4.000 398.440 ;
    END
  END i_dout0_1[6]
  PIN i_dout0_1[7]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 786.690 0.000 786.970 4.000 ;
    END
  END i_dout0_1[7]
  PIN i_dout0_1[8]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 806.010 0.000 806.290 4.000 ;
    END
  END i_dout0_1[8]
  PIN i_dout0_1[9]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 840.050 997.345 840.330 1001.345 ;
    END
  END i_dout0_1[9]
  PIN io_in[0]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 2.850 997.345 3.130 1001.345 ;
    END
  END io_in[0]
  PIN io_in[10]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 194.210 997.345 194.490 1001.345 ;
    END
  END io_in[10]
  PIN io_in[11]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 213.530 997.345 213.810 1001.345 ;
    END
  END io_in[11]
  PIN io_in[12]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 232.850 997.345 233.130 1001.345 ;
    END
  END io_in[12]
  PIN io_in[13]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 251.710 997.345 251.990 1001.345 ;
    END
  END io_in[13]
  PIN io_in[14]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 271.030 997.345 271.310 1001.345 ;
    END
  END io_in[14]
  PIN io_in[15]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 290.350 997.345 290.630 1001.345 ;
    END
  END io_in[15]
  PIN io_in[16]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 309.670 997.345 309.950 1001.345 ;
    END
  END io_in[16]
  PIN io_in[17]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 328.530 997.345 328.810 1001.345 ;
    END
  END io_in[17]
  PIN io_in[18]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 347.850 997.345 348.130 1001.345 ;
    END
  END io_in[18]
  PIN io_in[19]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 367.170 997.345 367.450 1001.345 ;
    END
  END io_in[19]
  PIN io_in[1]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 21.710 997.345 21.990 1001.345 ;
    END
  END io_in[1]
  PIN io_in[20]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 386.030 997.345 386.310 1001.345 ;
    END
  END io_in[20]
  PIN io_in[21]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 405.350 997.345 405.630 1001.345 ;
    END
  END io_in[21]
  PIN io_in[22]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 424.670 997.345 424.950 1001.345 ;
    END
  END io_in[22]
  PIN io_in[23]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 443.530 997.345 443.810 1001.345 ;
    END
  END io_in[23]
  PIN io_in[24]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 462.850 997.345 463.130 1001.345 ;
    END
  END io_in[24]
  PIN io_in[25]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 482.170 997.345 482.450 1001.345 ;
    END
  END io_in[25]
  PIN io_in[26]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 501.030 997.345 501.310 1001.345 ;
    END
  END io_in[26]
  PIN io_in[27]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 520.350 997.345 520.630 1001.345 ;
    END
  END io_in[27]
  PIN io_in[28]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 539.670 997.345 539.950 1001.345 ;
    END
  END io_in[28]
  PIN io_in[29]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 558.990 997.345 559.270 1001.345 ;
    END
  END io_in[29]
  PIN io_in[2]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 41.030 997.345 41.310 1001.345 ;
    END
  END io_in[2]
  PIN io_in[30]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 577.850 997.345 578.130 1001.345 ;
    END
  END io_in[30]
  PIN io_in[31]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 597.170 997.345 597.450 1001.345 ;
    END
  END io_in[31]
  PIN io_in[32]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 616.490 997.345 616.770 1001.345 ;
    END
  END io_in[32]
  PIN io_in[33]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 635.350 997.345 635.630 1001.345 ;
    END
  END io_in[33]
  PIN io_in[34]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 654.670 997.345 654.950 1001.345 ;
    END
  END io_in[34]
  PIN io_in[35]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 673.990 997.345 674.270 1001.345 ;
    END
  END io_in[35]
  PIN io_in[36]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 692.850 997.345 693.130 1001.345 ;
    END
  END io_in[36]
  PIN io_in[37]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 712.170 997.345 712.450 1001.345 ;
    END
  END io_in[37]
  PIN io_in[3]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 60.350 997.345 60.630 1001.345 ;
    END
  END io_in[3]
  PIN io_in[4]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 79.210 997.345 79.490 1001.345 ;
    END
  END io_in[4]
  PIN io_in[5]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 98.530 997.345 98.810 1001.345 ;
    END
  END io_in[5]
  PIN io_in[6]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 117.850 997.345 118.130 1001.345 ;
    END
  END io_in[6]
  PIN io_in[7]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 136.710 997.345 136.990 1001.345 ;
    END
  END io_in[7]
  PIN io_in[8]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 156.030 997.345 156.310 1001.345 ;
    END
  END io_in[8]
  PIN io_in[9]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 175.350 997.345 175.630 1001.345 ;
    END
  END io_in[9]
  PIN io_oeb[0]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 8.830 997.345 9.110 1001.345 ;
    END
  END io_oeb[0]
  PIN io_oeb[10]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 200.650 997.345 200.930 1001.345 ;
    END
  END io_oeb[10]
  PIN io_oeb[11]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 219.970 997.345 220.250 1001.345 ;
    END
  END io_oeb[11]
  PIN io_oeb[12]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 239.290 997.345 239.570 1001.345 ;
    END
  END io_oeb[12]
  PIN io_oeb[13]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 258.150 997.345 258.430 1001.345 ;
    END
  END io_oeb[13]
  PIN io_oeb[14]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 277.470 997.345 277.750 1001.345 ;
    END
  END io_oeb[14]
  PIN io_oeb[15]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 296.790 997.345 297.070 1001.345 ;
    END
  END io_oeb[15]
  PIN io_oeb[16]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 315.650 997.345 315.930 1001.345 ;
    END
  END io_oeb[16]
  PIN io_oeb[17]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 334.970 997.345 335.250 1001.345 ;
    END
  END io_oeb[17]
  PIN io_oeb[18]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 354.290 997.345 354.570 1001.345 ;
    END
  END io_oeb[18]
  PIN io_oeb[19]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 373.610 997.345 373.890 1001.345 ;
    END
  END io_oeb[19]
  PIN io_oeb[1]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 28.150 997.345 28.430 1001.345 ;
    END
  END io_oeb[1]
  PIN io_oeb[20]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 392.470 997.345 392.750 1001.345 ;
    END
  END io_oeb[20]
  PIN io_oeb[21]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 411.790 997.345 412.070 1001.345 ;
    END
  END io_oeb[21]
  PIN io_oeb[22]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 431.110 997.345 431.390 1001.345 ;
    END
  END io_oeb[22]
  PIN io_oeb[23]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 449.970 997.345 450.250 1001.345 ;
    END
  END io_oeb[23]
  PIN io_oeb[24]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 469.290 997.345 469.570 1001.345 ;
    END
  END io_oeb[24]
  PIN io_oeb[25]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 488.610 997.345 488.890 1001.345 ;
    END
  END io_oeb[25]
  PIN io_oeb[26]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 507.470 997.345 507.750 1001.345 ;
    END
  END io_oeb[26]
  PIN io_oeb[27]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 526.790 997.345 527.070 1001.345 ;
    END
  END io_oeb[27]
  PIN io_oeb[28]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 546.110 997.345 546.390 1001.345 ;
    END
  END io_oeb[28]
  PIN io_oeb[29]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 564.970 997.345 565.250 1001.345 ;
    END
  END io_oeb[29]
  PIN io_oeb[2]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 47.470 997.345 47.750 1001.345 ;
    END
  END io_oeb[2]
  PIN io_oeb[30]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 584.290 997.345 584.570 1001.345 ;
    END
  END io_oeb[30]
  PIN io_oeb[31]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 603.610 997.345 603.890 1001.345 ;
    END
  END io_oeb[31]
  PIN io_oeb[32]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 622.470 997.345 622.750 1001.345 ;
    END
  END io_oeb[32]
  PIN io_oeb[33]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 641.790 997.345 642.070 1001.345 ;
    END
  END io_oeb[33]
  PIN io_oeb[34]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 661.110 997.345 661.390 1001.345 ;
    END
  END io_oeb[34]
  PIN io_oeb[35]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 680.430 997.345 680.710 1001.345 ;
    END
  END io_oeb[35]
  PIN io_oeb[36]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 699.290 997.345 699.570 1001.345 ;
    END
  END io_oeb[36]
  PIN io_oeb[37]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 718.610 997.345 718.890 1001.345 ;
    END
  END io_oeb[37]
  PIN io_oeb[3]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 66.330 997.345 66.610 1001.345 ;
    END
  END io_oeb[3]
  PIN io_oeb[4]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 85.650 997.345 85.930 1001.345 ;
    END
  END io_oeb[4]
  PIN io_oeb[5]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 104.970 997.345 105.250 1001.345 ;
    END
  END io_oeb[5]
  PIN io_oeb[6]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 124.290 997.345 124.570 1001.345 ;
    END
  END io_oeb[6]
  PIN io_oeb[7]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 143.150 997.345 143.430 1001.345 ;
    END
  END io_oeb[7]
  PIN io_oeb[8]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 162.470 997.345 162.750 1001.345 ;
    END
  END io_oeb[8]
  PIN io_oeb[9]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 181.790 997.345 182.070 1001.345 ;
    END
  END io_oeb[9]
  PIN io_out[0]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 15.270 997.345 15.550 1001.345 ;
    END
  END io_out[0]
  PIN io_out[10]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 207.090 997.345 207.370 1001.345 ;
    END
  END io_out[10]
  PIN io_out[11]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 226.410 997.345 226.690 1001.345 ;
    END
  END io_out[11]
  PIN io_out[12]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 245.730 997.345 246.010 1001.345 ;
    END
  END io_out[12]
  PIN io_out[13]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 264.590 997.345 264.870 1001.345 ;
    END
  END io_out[13]
  PIN io_out[14]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 283.910 997.345 284.190 1001.345 ;
    END
  END io_out[14]
  PIN io_out[15]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 303.230 997.345 303.510 1001.345 ;
    END
  END io_out[15]
  PIN io_out[16]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 322.090 997.345 322.370 1001.345 ;
    END
  END io_out[16]
  PIN io_out[17]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 341.410 997.345 341.690 1001.345 ;
    END
  END io_out[17]
  PIN io_out[18]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 360.730 997.345 361.010 1001.345 ;
    END
  END io_out[18]
  PIN io_out[19]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 379.590 997.345 379.870 1001.345 ;
    END
  END io_out[19]
  PIN io_out[1]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 34.590 997.345 34.870 1001.345 ;
    END
  END io_out[1]
  PIN io_out[20]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 398.910 997.345 399.190 1001.345 ;
    END
  END io_out[20]
  PIN io_out[21]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 418.230 997.345 418.510 1001.345 ;
    END
  END io_out[21]
  PIN io_out[22]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 437.090 997.345 437.370 1001.345 ;
    END
  END io_out[22]
  PIN io_out[23]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 456.410 997.345 456.690 1001.345 ;
    END
  END io_out[23]
  PIN io_out[24]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 475.730 997.345 476.010 1001.345 ;
    END
  END io_out[24]
  PIN io_out[25]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 495.050 997.345 495.330 1001.345 ;
    END
  END io_out[25]
  PIN io_out[26]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 513.910 997.345 514.190 1001.345 ;
    END
  END io_out[26]
  PIN io_out[27]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 533.230 997.345 533.510 1001.345 ;
    END
  END io_out[27]
  PIN io_out[28]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 552.550 997.345 552.830 1001.345 ;
    END
  END io_out[28]
  PIN io_out[29]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 571.410 997.345 571.690 1001.345 ;
    END
  END io_out[29]
  PIN io_out[2]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 53.910 997.345 54.190 1001.345 ;
    END
  END io_out[2]
  PIN io_out[30]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 590.730 997.345 591.010 1001.345 ;
    END
  END io_out[30]
  PIN io_out[31]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 610.050 997.345 610.330 1001.345 ;
    END
  END io_out[31]
  PIN io_out[32]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 628.910 997.345 629.190 1001.345 ;
    END
  END io_out[32]
  PIN io_out[33]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 648.230 997.345 648.510 1001.345 ;
    END
  END io_out[33]
  PIN io_out[34]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 667.550 997.345 667.830 1001.345 ;
    END
  END io_out[34]
  PIN io_out[35]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 686.410 997.345 686.690 1001.345 ;
    END
  END io_out[35]
  PIN io_out[36]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 705.730 997.345 706.010 1001.345 ;
    END
  END io_out[36]
  PIN io_out[37]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 725.050 997.345 725.330 1001.345 ;
    END
  END io_out[37]
  PIN io_out[3]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 72.770 997.345 73.050 1001.345 ;
    END
  END io_out[3]
  PIN io_out[4]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 92.090 997.345 92.370 1001.345 ;
    END
  END io_out[4]
  PIN io_out[5]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 111.410 997.345 111.690 1001.345 ;
    END
  END io_out[5]
  PIN io_out[6]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 130.270 997.345 130.550 1001.345 ;
    END
  END io_out[6]
  PIN io_out[7]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 149.590 997.345 149.870 1001.345 ;
    END
  END io_out[7]
  PIN io_out[8]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 168.910 997.345 169.190 1001.345 ;
    END
  END io_out[8]
  PIN io_out[9]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 188.230 997.345 188.510 1001.345 ;
    END
  END io_out[9]
  PIN irq[0]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 689.630 0.000 689.910 4.000 ;
    END
  END irq[0]
  PIN irq[1]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 696.070 0.000 696.350 4.000 ;
    END
  END irq[1]
  PIN irq[2]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 702.510 0.000 702.790 4.000 ;
    END
  END irq[2]
  PIN o_csb0
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 10.920 4.000 11.520 ;
    END
  END o_csb0
  PIN o_csb0_1
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 986.625 47.640 990.625 48.240 ;
    END
  END o_csb0_1
  PIN o_din0[0]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 737.930 997.345 738.210 1001.345 ;
    END
  END o_din0[0]
  PIN o_din0[10]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 865.810 997.345 866.090 1001.345 ;
    END
  END o_din0[10]
  PIN o_din0[11]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 986.625 467.880 990.625 468.480 ;
    END
  END o_din0[11]
  PIN o_din0[12]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 857.990 0.000 858.270 4.000 ;
    END
  END o_din0[12]
  PIN o_din0[13]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 556.960 4.000 557.560 ;
    END
  END o_din0[13]
  PIN o_din0[14]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 870.870 0.000 871.150 4.000 ;
    END
  END o_din0[14]
  PIN o_din0[15]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 986.625 597.080 990.625 597.680 ;
    END
  END o_din0[15]
  PIN o_din0[16]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 986.625 629.040 990.625 629.640 ;
    END
  END o_din0[16]
  PIN o_din0[17]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 670.520 4.000 671.120 ;
    END
  END o_din0[17]
  PIN o_din0[18]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 716.080 4.000 716.680 ;
    END
  END o_din0[18]
  PIN o_din0[19]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 761.640 4.000 762.240 ;
    END
  END o_din0[19]
  PIN o_din0[1]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 750.350 997.345 750.630 1001.345 ;
    END
  END o_din0[1]
  PIN o_din0[20]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 784.760 4.000 785.360 ;
    END
  END o_din0[20]
  PIN o_din0[21]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 830.320 4.000 830.920 ;
    END
  END o_din0[21]
  PIN o_din0[22]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 986.625 822.840 990.625 823.440 ;
    END
  END o_din0[22]
  PIN o_din0[23]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 929.750 997.345 930.030 1001.345 ;
    END
  END o_din0[23]
  PIN o_din0[24]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 942.170 997.345 942.450 1001.345 ;
    END
  END o_din0[24]
  PIN o_din0[25]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 961.490 997.345 961.770 1001.345 ;
    END
  END o_din0[25]
  PIN o_din0[26]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 967.000 4.000 967.600 ;
    END
  END o_din0[26]
  PIN o_din0[27]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 929.290 0.000 929.570 4.000 ;
    END
  END o_din0[27]
  PIN o_din0[28]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 989.440 4.000 990.040 ;
    END
  END o_din0[28]
  PIN o_din0[29]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 986.625 952.040 990.625 952.640 ;
    END
  END o_din0[29]
  PIN o_din0[2]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 728.270 0.000 728.550 4.000 ;
    END
  END o_din0[2]
  PIN o_din0[30]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 974.370 0.000 974.650 4.000 ;
    END
  END o_din0[30]
  PIN o_din0[31]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 987.250 0.000 987.530 4.000 ;
    END
  END o_din0[31]
  PIN o_din0[3]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 986.625 274.080 990.625 274.680 ;
    END
  END o_din0[3]
  PIN o_din0[4]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 329.160 4.000 329.760 ;
    END
  END o_din0[4]
  PIN o_din0[5]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 352.280 4.000 352.880 ;
    END
  END o_din0[5]
  PIN o_din0[6]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 814.290 997.345 814.570 1001.345 ;
    END
  END o_din0[6]
  PIN o_din0[7]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 420.280 4.000 420.880 ;
    END
  END o_din0[7]
  PIN o_din0[8]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 465.840 4.000 466.440 ;
    END
  END o_din0[8]
  PIN o_din0[9]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 812.450 0.000 812.730 4.000 ;
    END
  END o_din0[9]
  PIN o_din0_1[0]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 744.370 997.345 744.650 1001.345 ;
    END
  END o_din0_1[0]
  PIN o_din0_1[10]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 859.370 997.345 859.650 1001.345 ;
    END
  END o_din0_1[10]
  PIN o_din0_1[11]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 986.625 435.240 990.625 435.840 ;
    END
  END o_din0_1[11]
  PIN o_din0_1[12]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 851.550 0.000 851.830 4.000 ;
    END
  END o_din0_1[12]
  PIN o_din0_1[13]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 871.790 997.345 872.070 1001.345 ;
    END
  END o_din0_1[13]
  PIN o_din0_1[14]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 864.430 0.000 864.710 4.000 ;
    END
  END o_din0_1[14]
  PIN o_din0_1[15]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 986.625 564.440 990.625 565.040 ;
    END
  END o_din0_1[15]
  PIN o_din0_1[16]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 891.110 997.345 891.390 1001.345 ;
    END
  END o_din0_1[16]
  PIN o_din0_1[17]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 883.750 0.000 884.030 4.000 ;
    END
  END o_din0_1[17]
  PIN o_din0_1[18]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 693.640 4.000 694.240 ;
    END
  END o_din0_1[18]
  PIN o_din0_1[19]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 986.625 693.640 990.625 694.240 ;
    END
  END o_din0_1[19]
  PIN o_din0_1[1]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 986.625 176.840 990.625 177.440 ;
    END
  END o_din0_1[1]
  PIN o_din0_1[20]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 910.430 997.345 910.710 1001.345 ;
    END
  END o_din0_1[20]
  PIN o_din0_1[21]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 986.625 758.240 990.625 758.840 ;
    END
  END o_din0_1[21]
  PIN o_din0_1[22]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 986.625 790.880 990.625 791.480 ;
    END
  END o_din0_1[22]
  PIN o_din0_1[23]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 986.625 855.480 990.625 856.080 ;
    END
  END o_din0_1[23]
  PIN o_din0_1[24]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 935.730 997.345 936.010 1001.345 ;
    END
  END o_din0_1[24]
  PIN o_din0_1[25]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 955.050 997.345 955.330 1001.345 ;
    END
  END o_din0_1[25]
  PIN o_din0_1[26]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 909.510 0.000 909.790 4.000 ;
    END
  END o_din0_1[26]
  PIN o_din0_1[27]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 986.625 887.440 990.625 888.040 ;
    END
  END o_din0_1[27]
  PIN o_din0_1[28]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 942.170 0.000 942.450 4.000 ;
    END
  END o_din0_1[28]
  PIN o_din0_1[29]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 948.610 0.000 948.890 4.000 ;
    END
  END o_din0_1[29]
  PIN o_din0_1[2]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 986.625 241.440 990.625 242.040 ;
    END
  END o_din0_1[2]
  PIN o_din0_1[30]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 967.930 0.000 968.210 4.000 ;
    END
  END o_din0_1[30]
  PIN o_din0_1[31]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 987.250 997.345 987.530 1001.345 ;
    END
  END o_din0_1[31]
  PIN o_din0_1[3]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 769.670 997.345 769.950 1001.345 ;
    END
  END o_din0_1[3]
  PIN o_din0_1[4]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 776.110 997.345 776.390 1001.345 ;
    END
  END o_din0_1[4]
  PIN o_din0_1[5]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 801.870 997.345 802.150 1001.345 ;
    END
  END o_din0_1[5]
  PIN o_din0_1[6]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 807.850 997.345 808.130 1001.345 ;
    END
  END o_din0_1[6]
  PIN o_din0_1[7]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 793.130 0.000 793.410 4.000 ;
    END
  END o_din0_1[7]
  PIN o_din0_1[8]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 986.625 403.280 990.625 403.880 ;
    END
  END o_din0_1[8]
  PIN o_din0_1[9]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 846.490 997.345 846.770 1001.345 ;
    END
  END o_din0_1[9]
  PIN o_waddr0[0]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 78.920 4.000 79.520 ;
    END
  END o_waddr0[0]
  PIN o_waddr0[1]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 721.830 0.000 722.110 4.000 ;
    END
  END o_waddr0[1]
  PIN o_waddr0[2]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 763.230 997.345 763.510 1001.345 ;
    END
  END o_waddr0[2]
  PIN o_waddr0[3]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 754.490 0.000 754.770 4.000 ;
    END
  END o_waddr0[3]
  PIN o_waddr0[4]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 788.990 997.345 789.270 1001.345 ;
    END
  END o_waddr0[4]
  PIN o_waddr0[5]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 773.810 0.000 774.090 4.000 ;
    END
  END o_waddr0[5]
  PIN o_waddr0[6]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 986.625 370.640 990.625 371.240 ;
    END
  END o_waddr0[6]
  PIN o_waddr0[7]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 799.570 0.000 799.850 4.000 ;
    END
  END o_waddr0[7]
  PIN o_waddr0[8]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 488.960 4.000 489.560 ;
    END
  END o_waddr0[8]
  PIN o_waddr0_1[0]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 101.360 4.000 101.960 ;
    END
  END o_waddr0_1[0]
  PIN o_waddr0_1[1]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 715.390 0.000 715.670 4.000 ;
    END
  END o_waddr0_1[1]
  PIN o_waddr0_1[2]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 756.790 997.345 757.070 1001.345 ;
    END
  END o_waddr0_1[2]
  PIN o_waddr0_1[3]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 261.160 4.000 261.760 ;
    END
  END o_waddr0_1[3]
  PIN o_waddr0_1[4]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 782.550 997.345 782.830 1001.345 ;
    END
  END o_waddr0_1[4]
  PIN o_waddr0_1[5]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 374.720 4.000 375.320 ;
    END
  END o_waddr0_1[5]
  PIN o_waddr0_1[6]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 780.250 0.000 780.530 4.000 ;
    END
  END o_waddr0_1[6]
  PIN o_waddr0_1[7]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 827.170 997.345 827.450 1001.345 ;
    END
  END o_waddr0_1[7]
  PIN o_waddr0_1[8]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 833.610 997.345 833.890 1001.345 ;
    END
  END o_waddr0_1[8]
  PIN o_web0
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 33.360 4.000 33.960 ;
    END
  END o_web0
  PIN o_web0_1
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 986.625 80.280 990.625 80.880 ;
    END
  END o_web0_1
  PIN o_wmask0[0]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 708.950 0.000 709.230 4.000 ;
    END
  END o_wmask0[0]
  PIN o_wmask0[1]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 192.480 4.000 193.080 ;
    END
  END o_wmask0[1]
  PIN o_wmask0[2]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 741.150 0.000 741.430 4.000 ;
    END
  END o_wmask0[2]
  PIN o_wmask0[3]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 283.600 4.000 284.200 ;
    END
  END o_wmask0[3]
  PIN o_wmask0_1[0]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 124.480 4.000 125.080 ;
    END
  END o_wmask0_1[0]
  PIN o_wmask0_1[1]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 170.040 4.000 170.640 ;
    END
  END o_wmask0_1[1]
  PIN o_wmask0_1[2]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 734.710 0.000 734.990 4.000 ;
    END
  END o_wmask0_1[2]
  PIN o_wmask0_1[3]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 760.930 0.000 761.210 4.000 ;
    END
  END o_wmask0_1[3]
  PIN rst_i
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 986.625 112.240 990.625 112.840 ;
    END
  END rst_i
  PIN vccd1
    DIRECTION INPUT ;
    USE POWER ;
    PORT
      LAYER met4 ;
        RECT 21.040 10.640 22.640 990.320 ;
    END
    PORT
      LAYER met4 ;
        RECT 174.640 10.640 176.240 990.320 ;
    END
    PORT
      LAYER met4 ;
        RECT 328.240 10.640 329.840 990.320 ;
    END
    PORT
      LAYER met4 ;
        RECT 481.840 10.640 483.440 990.320 ;
    END
    PORT
      LAYER met4 ;
        RECT 635.440 10.640 637.040 990.320 ;
    END
    PORT
      LAYER met4 ;
        RECT 789.040 10.640 790.640 990.320 ;
    END
    PORT
      LAYER met4 ;
        RECT 942.640 10.640 944.240 990.320 ;
    END
  END vccd1
  PIN vssd1
    DIRECTION INPUT ;
    USE GROUND ;
    PORT
      LAYER met4 ;
        RECT 97.840 10.640 99.440 990.320 ;
    END
    PORT
      LAYER met4 ;
        RECT 251.440 10.640 253.040 990.320 ;
    END
    PORT
      LAYER met4 ;
        RECT 405.040 10.640 406.640 990.320 ;
    END
    PORT
      LAYER met4 ;
        RECT 558.640 10.640 560.240 990.320 ;
    END
    PORT
      LAYER met4 ;
        RECT 712.240 10.640 713.840 990.320 ;
    END
    PORT
      LAYER met4 ;
        RECT 865.840 10.640 867.440 990.320 ;
    END
  END vssd1
  PIN wb_clk_i
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 3.310 0.000 3.590 4.000 ;
    END
  END wb_clk_i
  PIN wb_rst_i
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 9.750 0.000 10.030 4.000 ;
    END
  END wb_rst_i
  PIN wbs_ack_o
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 16.190 0.000 16.470 4.000 ;
    END
  END wbs_ack_o
  PIN wbs_adr_i[0]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 41.950 0.000 42.230 4.000 ;
    END
  END wbs_adr_i[0]
  PIN wbs_adr_i[10]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 262.290 0.000 262.570 4.000 ;
    END
  END wbs_adr_i[10]
  PIN wbs_adr_i[11]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 281.610 0.000 281.890 4.000 ;
    END
  END wbs_adr_i[11]
  PIN wbs_adr_i[12]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 300.930 0.000 301.210 4.000 ;
    END
  END wbs_adr_i[12]
  PIN wbs_adr_i[13]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 320.250 0.000 320.530 4.000 ;
    END
  END wbs_adr_i[13]
  PIN wbs_adr_i[14]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 340.030 0.000 340.310 4.000 ;
    END
  END wbs_adr_i[14]
  PIN wbs_adr_i[15]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 359.350 0.000 359.630 4.000 ;
    END
  END wbs_adr_i[15]
  PIN wbs_adr_i[16]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 378.670 0.000 378.950 4.000 ;
    END
  END wbs_adr_i[16]
  PIN wbs_adr_i[17]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 397.990 0.000 398.270 4.000 ;
    END
  END wbs_adr_i[17]
  PIN wbs_adr_i[18]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 417.770 0.000 418.050 4.000 ;
    END
  END wbs_adr_i[18]
  PIN wbs_adr_i[19]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 437.090 0.000 437.370 4.000 ;
    END
  END wbs_adr_i[19]
  PIN wbs_adr_i[1]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 67.710 0.000 67.990 4.000 ;
    END
  END wbs_adr_i[1]
  PIN wbs_adr_i[20]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 456.410 0.000 456.690 4.000 ;
    END
  END wbs_adr_i[20]
  PIN wbs_adr_i[21]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 475.730 0.000 476.010 4.000 ;
    END
  END wbs_adr_i[21]
  PIN wbs_adr_i[22]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 495.050 0.000 495.330 4.000 ;
    END
  END wbs_adr_i[22]
  PIN wbs_adr_i[23]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 514.830 0.000 515.110 4.000 ;
    END
  END wbs_adr_i[23]
  PIN wbs_adr_i[24]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 534.150 0.000 534.430 4.000 ;
    END
  END wbs_adr_i[24]
  PIN wbs_adr_i[25]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 553.470 0.000 553.750 4.000 ;
    END
  END wbs_adr_i[25]
  PIN wbs_adr_i[26]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 572.790 0.000 573.070 4.000 ;
    END
  END wbs_adr_i[26]
  PIN wbs_adr_i[27]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 592.570 0.000 592.850 4.000 ;
    END
  END wbs_adr_i[27]
  PIN wbs_adr_i[28]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 611.890 0.000 612.170 4.000 ;
    END
  END wbs_adr_i[28]
  PIN wbs_adr_i[29]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 631.210 0.000 631.490 4.000 ;
    END
  END wbs_adr_i[29]
  PIN wbs_adr_i[2]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 93.930 0.000 94.210 4.000 ;
    END
  END wbs_adr_i[2]
  PIN wbs_adr_i[30]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 650.530 0.000 650.810 4.000 ;
    END
  END wbs_adr_i[30]
  PIN wbs_adr_i[31]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 670.310 0.000 670.590 4.000 ;
    END
  END wbs_adr_i[31]
  PIN wbs_adr_i[3]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 119.690 0.000 119.970 4.000 ;
    END
  END wbs_adr_i[3]
  PIN wbs_adr_i[4]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 145.450 0.000 145.730 4.000 ;
    END
  END wbs_adr_i[4]
  PIN wbs_adr_i[5]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 164.770 0.000 165.050 4.000 ;
    END
  END wbs_adr_i[5]
  PIN wbs_adr_i[6]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 184.550 0.000 184.830 4.000 ;
    END
  END wbs_adr_i[6]
  PIN wbs_adr_i[7]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 203.870 0.000 204.150 4.000 ;
    END
  END wbs_adr_i[7]
  PIN wbs_adr_i[8]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 223.190 0.000 223.470 4.000 ;
    END
  END wbs_adr_i[8]
  PIN wbs_adr_i[9]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 242.510 0.000 242.790 4.000 ;
    END
  END wbs_adr_i[9]
  PIN wbs_cyc_i
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 22.630 0.000 22.910 4.000 ;
    END
  END wbs_cyc_i
  PIN wbs_dat_i[0]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 48.390 0.000 48.670 4.000 ;
    END
  END wbs_dat_i[0]
  PIN wbs_dat_i[10]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 268.730 0.000 269.010 4.000 ;
    END
  END wbs_dat_i[10]
  PIN wbs_dat_i[11]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 288.050 0.000 288.330 4.000 ;
    END
  END wbs_dat_i[11]
  PIN wbs_dat_i[12]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 307.370 0.000 307.650 4.000 ;
    END
  END wbs_dat_i[12]
  PIN wbs_dat_i[13]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 326.690 0.000 326.970 4.000 ;
    END
  END wbs_dat_i[13]
  PIN wbs_dat_i[14]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 346.470 0.000 346.750 4.000 ;
    END
  END wbs_dat_i[14]
  PIN wbs_dat_i[15]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 365.790 0.000 366.070 4.000 ;
    END
  END wbs_dat_i[15]
  PIN wbs_dat_i[16]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 385.110 0.000 385.390 4.000 ;
    END
  END wbs_dat_i[16]
  PIN wbs_dat_i[17]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 404.430 0.000 404.710 4.000 ;
    END
  END wbs_dat_i[17]
  PIN wbs_dat_i[18]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 424.210 0.000 424.490 4.000 ;
    END
  END wbs_dat_i[18]
  PIN wbs_dat_i[19]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 443.530 0.000 443.810 4.000 ;
    END
  END wbs_dat_i[19]
  PIN wbs_dat_i[1]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 74.150 0.000 74.430 4.000 ;
    END
  END wbs_dat_i[1]
  PIN wbs_dat_i[20]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 462.850 0.000 463.130 4.000 ;
    END
  END wbs_dat_i[20]
  PIN wbs_dat_i[21]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 482.170 0.000 482.450 4.000 ;
    END
  END wbs_dat_i[21]
  PIN wbs_dat_i[22]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 501.950 0.000 502.230 4.000 ;
    END
  END wbs_dat_i[22]
  PIN wbs_dat_i[23]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 521.270 0.000 521.550 4.000 ;
    END
  END wbs_dat_i[23]
  PIN wbs_dat_i[24]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 540.590 0.000 540.870 4.000 ;
    END
  END wbs_dat_i[24]
  PIN wbs_dat_i[25]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 559.910 0.000 560.190 4.000 ;
    END
  END wbs_dat_i[25]
  PIN wbs_dat_i[26]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 579.230 0.000 579.510 4.000 ;
    END
  END wbs_dat_i[26]
  PIN wbs_dat_i[27]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 599.010 0.000 599.290 4.000 ;
    END
  END wbs_dat_i[27]
  PIN wbs_dat_i[28]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 618.330 0.000 618.610 4.000 ;
    END
  END wbs_dat_i[28]
  PIN wbs_dat_i[29]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 637.650 0.000 637.930 4.000 ;
    END
  END wbs_dat_i[29]
  PIN wbs_dat_i[2]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 100.370 0.000 100.650 4.000 ;
    END
  END wbs_dat_i[2]
  PIN wbs_dat_i[30]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 656.970 0.000 657.250 4.000 ;
    END
  END wbs_dat_i[30]
  PIN wbs_dat_i[31]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 676.750 0.000 677.030 4.000 ;
    END
  END wbs_dat_i[31]
  PIN wbs_dat_i[3]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 126.130 0.000 126.410 4.000 ;
    END
  END wbs_dat_i[3]
  PIN wbs_dat_i[4]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 151.890 0.000 152.170 4.000 ;
    END
  END wbs_dat_i[4]
  PIN wbs_dat_i[5]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 171.670 0.000 171.950 4.000 ;
    END
  END wbs_dat_i[5]
  PIN wbs_dat_i[6]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 190.990 0.000 191.270 4.000 ;
    END
  END wbs_dat_i[6]
  PIN wbs_dat_i[7]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 210.310 0.000 210.590 4.000 ;
    END
  END wbs_dat_i[7]
  PIN wbs_dat_i[8]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 229.630 0.000 229.910 4.000 ;
    END
  END wbs_dat_i[8]
  PIN wbs_dat_i[9]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 248.950 0.000 249.230 4.000 ;
    END
  END wbs_dat_i[9]
  PIN wbs_dat_o[0]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 54.830 0.000 55.110 4.000 ;
    END
  END wbs_dat_o[0]
  PIN wbs_dat_o[10]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 275.170 0.000 275.450 4.000 ;
    END
  END wbs_dat_o[10]
  PIN wbs_dat_o[11]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 294.490 0.000 294.770 4.000 ;
    END
  END wbs_dat_o[11]
  PIN wbs_dat_o[12]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 313.810 0.000 314.090 4.000 ;
    END
  END wbs_dat_o[12]
  PIN wbs_dat_o[13]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 333.590 0.000 333.870 4.000 ;
    END
  END wbs_dat_o[13]
  PIN wbs_dat_o[14]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 352.910 0.000 353.190 4.000 ;
    END
  END wbs_dat_o[14]
  PIN wbs_dat_o[15]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 372.230 0.000 372.510 4.000 ;
    END
  END wbs_dat_o[15]
  PIN wbs_dat_o[16]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 391.550 0.000 391.830 4.000 ;
    END
  END wbs_dat_o[16]
  PIN wbs_dat_o[17]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 410.870 0.000 411.150 4.000 ;
    END
  END wbs_dat_o[17]
  PIN wbs_dat_o[18]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 430.650 0.000 430.930 4.000 ;
    END
  END wbs_dat_o[18]
  PIN wbs_dat_o[19]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 449.970 0.000 450.250 4.000 ;
    END
  END wbs_dat_o[19]
  PIN wbs_dat_o[1]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 80.590 0.000 80.870 4.000 ;
    END
  END wbs_dat_o[1]
  PIN wbs_dat_o[20]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 469.290 0.000 469.570 4.000 ;
    END
  END wbs_dat_o[20]
  PIN wbs_dat_o[21]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 488.610 0.000 488.890 4.000 ;
    END
  END wbs_dat_o[21]
  PIN wbs_dat_o[22]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 508.390 0.000 508.670 4.000 ;
    END
  END wbs_dat_o[22]
  PIN wbs_dat_o[23]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 527.710 0.000 527.990 4.000 ;
    END
  END wbs_dat_o[23]
  PIN wbs_dat_o[24]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 547.030 0.000 547.310 4.000 ;
    END
  END wbs_dat_o[24]
  PIN wbs_dat_o[25]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 566.350 0.000 566.630 4.000 ;
    END
  END wbs_dat_o[25]
  PIN wbs_dat_o[26]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 586.130 0.000 586.410 4.000 ;
    END
  END wbs_dat_o[26]
  PIN wbs_dat_o[27]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 605.450 0.000 605.730 4.000 ;
    END
  END wbs_dat_o[27]
  PIN wbs_dat_o[28]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 624.770 0.000 625.050 4.000 ;
    END
  END wbs_dat_o[28]
  PIN wbs_dat_o[29]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 644.090 0.000 644.370 4.000 ;
    END
  END wbs_dat_o[29]
  PIN wbs_dat_o[2]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 106.810 0.000 107.090 4.000 ;
    END
  END wbs_dat_o[2]
  PIN wbs_dat_o[30]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 663.870 0.000 664.150 4.000 ;
    END
  END wbs_dat_o[30]
  PIN wbs_dat_o[31]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 683.190 0.000 683.470 4.000 ;
    END
  END wbs_dat_o[31]
  PIN wbs_dat_o[3]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 132.570 0.000 132.850 4.000 ;
    END
  END wbs_dat_o[3]
  PIN wbs_dat_o[4]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 158.330 0.000 158.610 4.000 ;
    END
  END wbs_dat_o[4]
  PIN wbs_dat_o[5]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 178.110 0.000 178.390 4.000 ;
    END
  END wbs_dat_o[5]
  PIN wbs_dat_o[6]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 197.430 0.000 197.710 4.000 ;
    END
  END wbs_dat_o[6]
  PIN wbs_dat_o[7]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 216.750 0.000 217.030 4.000 ;
    END
  END wbs_dat_o[7]
  PIN wbs_dat_o[8]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 236.070 0.000 236.350 4.000 ;
    END
  END wbs_dat_o[8]
  PIN wbs_dat_o[9]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 255.850 0.000 256.130 4.000 ;
    END
  END wbs_dat_o[9]
  PIN wbs_sel_i[0]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 61.270 0.000 61.550 4.000 ;
    END
  END wbs_sel_i[0]
  PIN wbs_sel_i[1]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 87.490 0.000 87.770 4.000 ;
    END
  END wbs_sel_i[1]
  PIN wbs_sel_i[2]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 113.250 0.000 113.530 4.000 ;
    END
  END wbs_sel_i[2]
  PIN wbs_sel_i[3]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 139.010 0.000 139.290 4.000 ;
    END
  END wbs_sel_i[3]
  PIN wbs_stb_i
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 29.070 0.000 29.350 4.000 ;
    END
  END wbs_stb_i
  PIN wbs_we_i
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 35.510 0.000 35.790 4.000 ;
    END
  END wbs_we_i
  OBS
      LAYER li1 ;
        RECT 5.520 10.795 987.015 990.165 ;
      LAYER met1 ;
        RECT 3.290 4.800 988.470 991.060 ;
      LAYER met2 ;
        RECT 3.410 997.065 8.550 997.345 ;
        RECT 9.390 997.065 14.990 997.345 ;
        RECT 15.830 997.065 21.430 997.345 ;
        RECT 22.270 997.065 27.870 997.345 ;
        RECT 28.710 997.065 34.310 997.345 ;
        RECT 35.150 997.065 40.750 997.345 ;
        RECT 41.590 997.065 47.190 997.345 ;
        RECT 48.030 997.065 53.630 997.345 ;
        RECT 54.470 997.065 60.070 997.345 ;
        RECT 60.910 997.065 66.050 997.345 ;
        RECT 66.890 997.065 72.490 997.345 ;
        RECT 73.330 997.065 78.930 997.345 ;
        RECT 79.770 997.065 85.370 997.345 ;
        RECT 86.210 997.065 91.810 997.345 ;
        RECT 92.650 997.065 98.250 997.345 ;
        RECT 99.090 997.065 104.690 997.345 ;
        RECT 105.530 997.065 111.130 997.345 ;
        RECT 111.970 997.065 117.570 997.345 ;
        RECT 118.410 997.065 124.010 997.345 ;
        RECT 124.850 997.065 129.990 997.345 ;
        RECT 130.830 997.065 136.430 997.345 ;
        RECT 137.270 997.065 142.870 997.345 ;
        RECT 143.710 997.065 149.310 997.345 ;
        RECT 150.150 997.065 155.750 997.345 ;
        RECT 156.590 997.065 162.190 997.345 ;
        RECT 163.030 997.065 168.630 997.345 ;
        RECT 169.470 997.065 175.070 997.345 ;
        RECT 175.910 997.065 181.510 997.345 ;
        RECT 182.350 997.065 187.950 997.345 ;
        RECT 188.790 997.065 193.930 997.345 ;
        RECT 194.770 997.065 200.370 997.345 ;
        RECT 201.210 997.065 206.810 997.345 ;
        RECT 207.650 997.065 213.250 997.345 ;
        RECT 214.090 997.065 219.690 997.345 ;
        RECT 220.530 997.065 226.130 997.345 ;
        RECT 226.970 997.065 232.570 997.345 ;
        RECT 233.410 997.065 239.010 997.345 ;
        RECT 239.850 997.065 245.450 997.345 ;
        RECT 246.290 997.065 251.430 997.345 ;
        RECT 252.270 997.065 257.870 997.345 ;
        RECT 258.710 997.065 264.310 997.345 ;
        RECT 265.150 997.065 270.750 997.345 ;
        RECT 271.590 997.065 277.190 997.345 ;
        RECT 278.030 997.065 283.630 997.345 ;
        RECT 284.470 997.065 290.070 997.345 ;
        RECT 290.910 997.065 296.510 997.345 ;
        RECT 297.350 997.065 302.950 997.345 ;
        RECT 303.790 997.065 309.390 997.345 ;
        RECT 310.230 997.065 315.370 997.345 ;
        RECT 316.210 997.065 321.810 997.345 ;
        RECT 322.650 997.065 328.250 997.345 ;
        RECT 329.090 997.065 334.690 997.345 ;
        RECT 335.530 997.065 341.130 997.345 ;
        RECT 341.970 997.065 347.570 997.345 ;
        RECT 348.410 997.065 354.010 997.345 ;
        RECT 354.850 997.065 360.450 997.345 ;
        RECT 361.290 997.065 366.890 997.345 ;
        RECT 367.730 997.065 373.330 997.345 ;
        RECT 374.170 997.065 379.310 997.345 ;
        RECT 380.150 997.065 385.750 997.345 ;
        RECT 386.590 997.065 392.190 997.345 ;
        RECT 393.030 997.065 398.630 997.345 ;
        RECT 399.470 997.065 405.070 997.345 ;
        RECT 405.910 997.065 411.510 997.345 ;
        RECT 412.350 997.065 417.950 997.345 ;
        RECT 418.790 997.065 424.390 997.345 ;
        RECT 425.230 997.065 430.830 997.345 ;
        RECT 431.670 997.065 436.810 997.345 ;
        RECT 437.650 997.065 443.250 997.345 ;
        RECT 444.090 997.065 449.690 997.345 ;
        RECT 450.530 997.065 456.130 997.345 ;
        RECT 456.970 997.065 462.570 997.345 ;
        RECT 463.410 997.065 469.010 997.345 ;
        RECT 469.850 997.065 475.450 997.345 ;
        RECT 476.290 997.065 481.890 997.345 ;
        RECT 482.730 997.065 488.330 997.345 ;
        RECT 489.170 997.065 494.770 997.345 ;
        RECT 495.610 997.065 500.750 997.345 ;
        RECT 501.590 997.065 507.190 997.345 ;
        RECT 508.030 997.065 513.630 997.345 ;
        RECT 514.470 997.065 520.070 997.345 ;
        RECT 520.910 997.065 526.510 997.345 ;
        RECT 527.350 997.065 532.950 997.345 ;
        RECT 533.790 997.065 539.390 997.345 ;
        RECT 540.230 997.065 545.830 997.345 ;
        RECT 546.670 997.065 552.270 997.345 ;
        RECT 553.110 997.065 558.710 997.345 ;
        RECT 559.550 997.065 564.690 997.345 ;
        RECT 565.530 997.065 571.130 997.345 ;
        RECT 571.970 997.065 577.570 997.345 ;
        RECT 578.410 997.065 584.010 997.345 ;
        RECT 584.850 997.065 590.450 997.345 ;
        RECT 591.290 997.065 596.890 997.345 ;
        RECT 597.730 997.065 603.330 997.345 ;
        RECT 604.170 997.065 609.770 997.345 ;
        RECT 610.610 997.065 616.210 997.345 ;
        RECT 617.050 997.065 622.190 997.345 ;
        RECT 623.030 997.065 628.630 997.345 ;
        RECT 629.470 997.065 635.070 997.345 ;
        RECT 635.910 997.065 641.510 997.345 ;
        RECT 642.350 997.065 647.950 997.345 ;
        RECT 648.790 997.065 654.390 997.345 ;
        RECT 655.230 997.065 660.830 997.345 ;
        RECT 661.670 997.065 667.270 997.345 ;
        RECT 668.110 997.065 673.710 997.345 ;
        RECT 674.550 997.065 680.150 997.345 ;
        RECT 680.990 997.065 686.130 997.345 ;
        RECT 686.970 997.065 692.570 997.345 ;
        RECT 693.410 997.065 699.010 997.345 ;
        RECT 699.850 997.065 705.450 997.345 ;
        RECT 706.290 997.065 711.890 997.345 ;
        RECT 712.730 997.065 718.330 997.345 ;
        RECT 719.170 997.065 724.770 997.345 ;
        RECT 725.610 997.065 731.210 997.345 ;
        RECT 732.050 997.065 737.650 997.345 ;
        RECT 738.490 997.065 744.090 997.345 ;
        RECT 744.930 997.065 750.070 997.345 ;
        RECT 750.910 997.065 756.510 997.345 ;
        RECT 757.350 997.065 762.950 997.345 ;
        RECT 763.790 997.065 769.390 997.345 ;
        RECT 770.230 997.065 775.830 997.345 ;
        RECT 776.670 997.065 782.270 997.345 ;
        RECT 783.110 997.065 788.710 997.345 ;
        RECT 789.550 997.065 795.150 997.345 ;
        RECT 795.990 997.065 801.590 997.345 ;
        RECT 802.430 997.065 807.570 997.345 ;
        RECT 808.410 997.065 814.010 997.345 ;
        RECT 814.850 997.065 820.450 997.345 ;
        RECT 821.290 997.065 826.890 997.345 ;
        RECT 827.730 997.065 833.330 997.345 ;
        RECT 834.170 997.065 839.770 997.345 ;
        RECT 840.610 997.065 846.210 997.345 ;
        RECT 847.050 997.065 852.650 997.345 ;
        RECT 853.490 997.065 859.090 997.345 ;
        RECT 859.930 997.065 865.530 997.345 ;
        RECT 866.370 997.065 871.510 997.345 ;
        RECT 872.350 997.065 877.950 997.345 ;
        RECT 878.790 997.065 884.390 997.345 ;
        RECT 885.230 997.065 890.830 997.345 ;
        RECT 891.670 997.065 897.270 997.345 ;
        RECT 898.110 997.065 903.710 997.345 ;
        RECT 904.550 997.065 910.150 997.345 ;
        RECT 910.990 997.065 916.590 997.345 ;
        RECT 917.430 997.065 923.030 997.345 ;
        RECT 923.870 997.065 929.470 997.345 ;
        RECT 930.310 997.065 935.450 997.345 ;
        RECT 936.290 997.065 941.890 997.345 ;
        RECT 942.730 997.065 948.330 997.345 ;
        RECT 949.170 997.065 954.770 997.345 ;
        RECT 955.610 997.065 961.210 997.345 ;
        RECT 962.050 997.065 967.650 997.345 ;
        RECT 968.490 997.065 974.090 997.345 ;
        RECT 974.930 997.065 980.530 997.345 ;
        RECT 981.370 997.065 986.970 997.345 ;
        RECT 987.810 997.065 988.450 997.345 ;
        RECT 3.320 4.280 988.450 997.065 ;
        RECT 3.870 3.670 9.470 4.280 ;
        RECT 10.310 3.670 15.910 4.280 ;
        RECT 16.750 3.670 22.350 4.280 ;
        RECT 23.190 3.670 28.790 4.280 ;
        RECT 29.630 3.670 35.230 4.280 ;
        RECT 36.070 3.670 41.670 4.280 ;
        RECT 42.510 3.670 48.110 4.280 ;
        RECT 48.950 3.670 54.550 4.280 ;
        RECT 55.390 3.670 60.990 4.280 ;
        RECT 61.830 3.670 67.430 4.280 ;
        RECT 68.270 3.670 73.870 4.280 ;
        RECT 74.710 3.670 80.310 4.280 ;
        RECT 81.150 3.670 87.210 4.280 ;
        RECT 88.050 3.670 93.650 4.280 ;
        RECT 94.490 3.670 100.090 4.280 ;
        RECT 100.930 3.670 106.530 4.280 ;
        RECT 107.370 3.670 112.970 4.280 ;
        RECT 113.810 3.670 119.410 4.280 ;
        RECT 120.250 3.670 125.850 4.280 ;
        RECT 126.690 3.670 132.290 4.280 ;
        RECT 133.130 3.670 138.730 4.280 ;
        RECT 139.570 3.670 145.170 4.280 ;
        RECT 146.010 3.670 151.610 4.280 ;
        RECT 152.450 3.670 158.050 4.280 ;
        RECT 158.890 3.670 164.490 4.280 ;
        RECT 165.330 3.670 171.390 4.280 ;
        RECT 172.230 3.670 177.830 4.280 ;
        RECT 178.670 3.670 184.270 4.280 ;
        RECT 185.110 3.670 190.710 4.280 ;
        RECT 191.550 3.670 197.150 4.280 ;
        RECT 197.990 3.670 203.590 4.280 ;
        RECT 204.430 3.670 210.030 4.280 ;
        RECT 210.870 3.670 216.470 4.280 ;
        RECT 217.310 3.670 222.910 4.280 ;
        RECT 223.750 3.670 229.350 4.280 ;
        RECT 230.190 3.670 235.790 4.280 ;
        RECT 236.630 3.670 242.230 4.280 ;
        RECT 243.070 3.670 248.670 4.280 ;
        RECT 249.510 3.670 255.570 4.280 ;
        RECT 256.410 3.670 262.010 4.280 ;
        RECT 262.850 3.670 268.450 4.280 ;
        RECT 269.290 3.670 274.890 4.280 ;
        RECT 275.730 3.670 281.330 4.280 ;
        RECT 282.170 3.670 287.770 4.280 ;
        RECT 288.610 3.670 294.210 4.280 ;
        RECT 295.050 3.670 300.650 4.280 ;
        RECT 301.490 3.670 307.090 4.280 ;
        RECT 307.930 3.670 313.530 4.280 ;
        RECT 314.370 3.670 319.970 4.280 ;
        RECT 320.810 3.670 326.410 4.280 ;
        RECT 327.250 3.670 333.310 4.280 ;
        RECT 334.150 3.670 339.750 4.280 ;
        RECT 340.590 3.670 346.190 4.280 ;
        RECT 347.030 3.670 352.630 4.280 ;
        RECT 353.470 3.670 359.070 4.280 ;
        RECT 359.910 3.670 365.510 4.280 ;
        RECT 366.350 3.670 371.950 4.280 ;
        RECT 372.790 3.670 378.390 4.280 ;
        RECT 379.230 3.670 384.830 4.280 ;
        RECT 385.670 3.670 391.270 4.280 ;
        RECT 392.110 3.670 397.710 4.280 ;
        RECT 398.550 3.670 404.150 4.280 ;
        RECT 404.990 3.670 410.590 4.280 ;
        RECT 411.430 3.670 417.490 4.280 ;
        RECT 418.330 3.670 423.930 4.280 ;
        RECT 424.770 3.670 430.370 4.280 ;
        RECT 431.210 3.670 436.810 4.280 ;
        RECT 437.650 3.670 443.250 4.280 ;
        RECT 444.090 3.670 449.690 4.280 ;
        RECT 450.530 3.670 456.130 4.280 ;
        RECT 456.970 3.670 462.570 4.280 ;
        RECT 463.410 3.670 469.010 4.280 ;
        RECT 469.850 3.670 475.450 4.280 ;
        RECT 476.290 3.670 481.890 4.280 ;
        RECT 482.730 3.670 488.330 4.280 ;
        RECT 489.170 3.670 494.770 4.280 ;
        RECT 495.610 3.670 501.670 4.280 ;
        RECT 502.510 3.670 508.110 4.280 ;
        RECT 508.950 3.670 514.550 4.280 ;
        RECT 515.390 3.670 520.990 4.280 ;
        RECT 521.830 3.670 527.430 4.280 ;
        RECT 528.270 3.670 533.870 4.280 ;
        RECT 534.710 3.670 540.310 4.280 ;
        RECT 541.150 3.670 546.750 4.280 ;
        RECT 547.590 3.670 553.190 4.280 ;
        RECT 554.030 3.670 559.630 4.280 ;
        RECT 560.470 3.670 566.070 4.280 ;
        RECT 566.910 3.670 572.510 4.280 ;
        RECT 573.350 3.670 578.950 4.280 ;
        RECT 579.790 3.670 585.850 4.280 ;
        RECT 586.690 3.670 592.290 4.280 ;
        RECT 593.130 3.670 598.730 4.280 ;
        RECT 599.570 3.670 605.170 4.280 ;
        RECT 606.010 3.670 611.610 4.280 ;
        RECT 612.450 3.670 618.050 4.280 ;
        RECT 618.890 3.670 624.490 4.280 ;
        RECT 625.330 3.670 630.930 4.280 ;
        RECT 631.770 3.670 637.370 4.280 ;
        RECT 638.210 3.670 643.810 4.280 ;
        RECT 644.650 3.670 650.250 4.280 ;
        RECT 651.090 3.670 656.690 4.280 ;
        RECT 657.530 3.670 663.590 4.280 ;
        RECT 664.430 3.670 670.030 4.280 ;
        RECT 670.870 3.670 676.470 4.280 ;
        RECT 677.310 3.670 682.910 4.280 ;
        RECT 683.750 3.670 689.350 4.280 ;
        RECT 690.190 3.670 695.790 4.280 ;
        RECT 696.630 3.670 702.230 4.280 ;
        RECT 703.070 3.670 708.670 4.280 ;
        RECT 709.510 3.670 715.110 4.280 ;
        RECT 715.950 3.670 721.550 4.280 ;
        RECT 722.390 3.670 727.990 4.280 ;
        RECT 728.830 3.670 734.430 4.280 ;
        RECT 735.270 3.670 740.870 4.280 ;
        RECT 741.710 3.670 747.770 4.280 ;
        RECT 748.610 3.670 754.210 4.280 ;
        RECT 755.050 3.670 760.650 4.280 ;
        RECT 761.490 3.670 767.090 4.280 ;
        RECT 767.930 3.670 773.530 4.280 ;
        RECT 774.370 3.670 779.970 4.280 ;
        RECT 780.810 3.670 786.410 4.280 ;
        RECT 787.250 3.670 792.850 4.280 ;
        RECT 793.690 3.670 799.290 4.280 ;
        RECT 800.130 3.670 805.730 4.280 ;
        RECT 806.570 3.670 812.170 4.280 ;
        RECT 813.010 3.670 818.610 4.280 ;
        RECT 819.450 3.670 825.050 4.280 ;
        RECT 825.890 3.670 831.950 4.280 ;
        RECT 832.790 3.670 838.390 4.280 ;
        RECT 839.230 3.670 844.830 4.280 ;
        RECT 845.670 3.670 851.270 4.280 ;
        RECT 852.110 3.670 857.710 4.280 ;
        RECT 858.550 3.670 864.150 4.280 ;
        RECT 864.990 3.670 870.590 4.280 ;
        RECT 871.430 3.670 877.030 4.280 ;
        RECT 877.870 3.670 883.470 4.280 ;
        RECT 884.310 3.670 889.910 4.280 ;
        RECT 890.750 3.670 896.350 4.280 ;
        RECT 897.190 3.670 902.790 4.280 ;
        RECT 903.630 3.670 909.230 4.280 ;
        RECT 910.070 3.670 916.130 4.280 ;
        RECT 916.970 3.670 922.570 4.280 ;
        RECT 923.410 3.670 929.010 4.280 ;
        RECT 929.850 3.670 935.450 4.280 ;
        RECT 936.290 3.670 941.890 4.280 ;
        RECT 942.730 3.670 948.330 4.280 ;
        RECT 949.170 3.670 954.770 4.280 ;
        RECT 955.610 3.670 961.210 4.280 ;
        RECT 962.050 3.670 967.650 4.280 ;
        RECT 968.490 3.670 974.090 4.280 ;
        RECT 974.930 3.670 980.530 4.280 ;
        RECT 981.370 3.670 986.970 4.280 ;
        RECT 987.810 3.670 988.450 4.280 ;
      LAYER met3 ;
        RECT 4.000 990.440 988.475 991.945 ;
        RECT 4.400 989.040 988.475 990.440 ;
        RECT 4.000 985.680 988.475 989.040 ;
        RECT 4.000 984.280 986.225 985.680 ;
        RECT 4.000 968.000 988.475 984.280 ;
        RECT 4.400 966.600 988.475 968.000 ;
        RECT 4.000 953.040 988.475 966.600 ;
        RECT 4.000 951.640 986.225 953.040 ;
        RECT 4.000 944.880 988.475 951.640 ;
        RECT 4.400 943.480 988.475 944.880 ;
        RECT 4.000 922.440 988.475 943.480 ;
        RECT 4.400 921.080 988.475 922.440 ;
        RECT 4.400 921.040 986.225 921.080 ;
        RECT 4.000 919.680 986.225 921.040 ;
        RECT 4.000 899.320 988.475 919.680 ;
        RECT 4.400 897.920 988.475 899.320 ;
        RECT 4.000 888.440 988.475 897.920 ;
        RECT 4.000 887.040 986.225 888.440 ;
        RECT 4.000 876.880 988.475 887.040 ;
        RECT 4.400 875.480 988.475 876.880 ;
        RECT 4.000 856.480 988.475 875.480 ;
        RECT 4.000 855.080 986.225 856.480 ;
        RECT 4.000 853.760 988.475 855.080 ;
        RECT 4.400 852.360 988.475 853.760 ;
        RECT 4.000 831.320 988.475 852.360 ;
        RECT 4.400 829.920 988.475 831.320 ;
        RECT 4.000 823.840 988.475 829.920 ;
        RECT 4.000 822.440 986.225 823.840 ;
        RECT 4.000 808.200 988.475 822.440 ;
        RECT 4.400 806.800 988.475 808.200 ;
        RECT 4.000 791.880 988.475 806.800 ;
        RECT 4.000 790.480 986.225 791.880 ;
        RECT 4.000 785.760 988.475 790.480 ;
        RECT 4.400 784.360 988.475 785.760 ;
        RECT 4.000 762.640 988.475 784.360 ;
        RECT 4.400 761.240 988.475 762.640 ;
        RECT 4.000 759.240 988.475 761.240 ;
        RECT 4.000 757.840 986.225 759.240 ;
        RECT 4.000 740.200 988.475 757.840 ;
        RECT 4.400 738.800 988.475 740.200 ;
        RECT 4.000 727.280 988.475 738.800 ;
        RECT 4.000 725.880 986.225 727.280 ;
        RECT 4.000 717.080 988.475 725.880 ;
        RECT 4.400 715.680 988.475 717.080 ;
        RECT 4.000 694.640 988.475 715.680 ;
        RECT 4.400 693.240 986.225 694.640 ;
        RECT 4.000 671.520 988.475 693.240 ;
        RECT 4.400 670.120 988.475 671.520 ;
        RECT 4.000 662.680 988.475 670.120 ;
        RECT 4.000 661.280 986.225 662.680 ;
        RECT 4.000 649.080 988.475 661.280 ;
        RECT 4.400 647.680 988.475 649.080 ;
        RECT 4.000 630.040 988.475 647.680 ;
        RECT 4.000 628.640 986.225 630.040 ;
        RECT 4.000 625.960 988.475 628.640 ;
        RECT 4.400 624.560 988.475 625.960 ;
        RECT 4.000 603.520 988.475 624.560 ;
        RECT 4.400 602.120 988.475 603.520 ;
        RECT 4.000 598.080 988.475 602.120 ;
        RECT 4.000 596.680 986.225 598.080 ;
        RECT 4.000 580.400 988.475 596.680 ;
        RECT 4.400 579.000 988.475 580.400 ;
        RECT 4.000 565.440 988.475 579.000 ;
        RECT 4.000 564.040 986.225 565.440 ;
        RECT 4.000 557.960 988.475 564.040 ;
        RECT 4.400 556.560 988.475 557.960 ;
        RECT 4.000 534.840 988.475 556.560 ;
        RECT 4.400 533.480 988.475 534.840 ;
        RECT 4.400 533.440 986.225 533.480 ;
        RECT 4.000 532.080 986.225 533.440 ;
        RECT 4.000 512.400 988.475 532.080 ;
        RECT 4.400 511.000 988.475 512.400 ;
        RECT 4.000 500.840 988.475 511.000 ;
        RECT 4.000 499.440 986.225 500.840 ;
        RECT 4.000 489.960 988.475 499.440 ;
        RECT 4.400 488.560 988.475 489.960 ;
        RECT 4.000 468.880 988.475 488.560 ;
        RECT 4.000 467.480 986.225 468.880 ;
        RECT 4.000 466.840 988.475 467.480 ;
        RECT 4.400 465.440 988.475 466.840 ;
        RECT 4.000 444.400 988.475 465.440 ;
        RECT 4.400 443.000 988.475 444.400 ;
        RECT 4.000 436.240 988.475 443.000 ;
        RECT 4.000 434.840 986.225 436.240 ;
        RECT 4.000 421.280 988.475 434.840 ;
        RECT 4.400 419.880 988.475 421.280 ;
        RECT 4.000 404.280 988.475 419.880 ;
        RECT 4.000 402.880 986.225 404.280 ;
        RECT 4.000 398.840 988.475 402.880 ;
        RECT 4.400 397.440 988.475 398.840 ;
        RECT 4.000 375.720 988.475 397.440 ;
        RECT 4.400 374.320 988.475 375.720 ;
        RECT 4.000 371.640 988.475 374.320 ;
        RECT 4.000 370.240 986.225 371.640 ;
        RECT 4.000 353.280 988.475 370.240 ;
        RECT 4.400 351.880 988.475 353.280 ;
        RECT 4.000 339.680 988.475 351.880 ;
        RECT 4.000 338.280 986.225 339.680 ;
        RECT 4.000 330.160 988.475 338.280 ;
        RECT 4.400 328.760 988.475 330.160 ;
        RECT 4.000 307.720 988.475 328.760 ;
        RECT 4.400 307.040 988.475 307.720 ;
        RECT 4.400 306.320 986.225 307.040 ;
        RECT 4.000 305.640 986.225 306.320 ;
        RECT 4.000 284.600 988.475 305.640 ;
        RECT 4.400 283.200 988.475 284.600 ;
        RECT 4.000 275.080 988.475 283.200 ;
        RECT 4.000 273.680 986.225 275.080 ;
        RECT 4.000 262.160 988.475 273.680 ;
        RECT 4.400 260.760 988.475 262.160 ;
        RECT 4.000 242.440 988.475 260.760 ;
        RECT 4.000 241.040 986.225 242.440 ;
        RECT 4.000 239.040 988.475 241.040 ;
        RECT 4.400 237.640 988.475 239.040 ;
        RECT 4.000 216.600 988.475 237.640 ;
        RECT 4.400 215.200 988.475 216.600 ;
        RECT 4.000 210.480 988.475 215.200 ;
        RECT 4.000 209.080 986.225 210.480 ;
        RECT 4.000 193.480 988.475 209.080 ;
        RECT 4.400 192.080 988.475 193.480 ;
        RECT 4.000 177.840 988.475 192.080 ;
        RECT 4.000 176.440 986.225 177.840 ;
        RECT 4.000 171.040 988.475 176.440 ;
        RECT 4.400 169.640 988.475 171.040 ;
        RECT 4.000 147.920 988.475 169.640 ;
        RECT 4.400 146.520 988.475 147.920 ;
        RECT 4.000 145.880 988.475 146.520 ;
        RECT 4.000 144.480 986.225 145.880 ;
        RECT 4.000 125.480 988.475 144.480 ;
        RECT 4.400 124.080 988.475 125.480 ;
        RECT 4.000 113.240 988.475 124.080 ;
        RECT 4.000 111.840 986.225 113.240 ;
        RECT 4.000 102.360 988.475 111.840 ;
        RECT 4.400 100.960 988.475 102.360 ;
        RECT 4.000 81.280 988.475 100.960 ;
        RECT 4.000 79.920 986.225 81.280 ;
        RECT 4.400 79.880 986.225 79.920 ;
        RECT 4.400 78.520 988.475 79.880 ;
        RECT 4.000 56.800 988.475 78.520 ;
        RECT 4.400 55.400 988.475 56.800 ;
        RECT 4.000 48.640 988.475 55.400 ;
        RECT 4.000 47.240 986.225 48.640 ;
        RECT 4.000 34.360 988.475 47.240 ;
        RECT 4.400 32.960 988.475 34.360 ;
        RECT 4.000 16.680 988.475 32.960 ;
        RECT 4.000 15.280 986.225 16.680 ;
        RECT 4.000 11.920 988.475 15.280 ;
        RECT 4.400 10.715 988.475 11.920 ;
      LAYER met4 ;
        RECT 54.575 990.720 977.665 991.945 ;
        RECT 54.575 14.455 97.440 990.720 ;
        RECT 99.840 14.455 174.240 990.720 ;
        RECT 176.640 14.455 251.040 990.720 ;
        RECT 253.440 14.455 327.840 990.720 ;
        RECT 330.240 14.455 404.640 990.720 ;
        RECT 407.040 14.455 481.440 990.720 ;
        RECT 483.840 14.455 558.240 990.720 ;
        RECT 560.640 14.455 635.040 990.720 ;
        RECT 637.440 14.455 711.840 990.720 ;
        RECT 714.240 14.455 788.640 990.720 ;
        RECT 791.040 14.455 865.440 990.720 ;
        RECT 867.840 14.455 942.240 990.720 ;
        RECT 944.640 14.455 977.665 990.720 ;
  END
END user_proj
END LIBRARY

